`timescale 1ns / 1ps

package Board_params;

    parameter NET_CLOCK_PERIOD = 3.1; // in ns
    parameter MAC_CLOCK_PERIOD = 3.1; // in ns

    parameter NET_DATA_WIDTH = 512;
  
endpackage
