/*

Copyright (c) 2014-2021 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall `timescale 1ns / 1ps `default_nettype none

/*
 * FPGA core logic
 */
module top (
    /*
     * Clock: 390.625 MHz
     * Synchronous reset
     */
    input wire clk,
    input wire rst,

    /*
     * GPIO
     */
    input  wire       btnu,
    input  wire       btnl,
    input  wire       btnd,
    input  wire       btnr,
    input  wire       btnc,
    input  wire [3:0] sw,
    output wire [7:0] led,

    /*
     * Ethernet: QSFP28
     */
    input  wire        xgmii_tx_clk,
    input  wire        xgmii_tx_rst,
    output wire [63:0] xgmii_txd,
    output wire [ 7:0] xgmii_txc,
    input  wire        xgmii_rx_clk,
    input  wire        xgmii_rx_rst,
    input  wire [63:0] xgmii_rxd,
    input  wire [ 7:0] xgmii_rxc
);


  wire [63:0] rx_axis_tdata;
  wire [7:0] rx_axis_tkeep;
  wire rx_axis_tvalid;
  wire rx_axis_tready;
  wire rx_axis_tlast;
  wire rx_axis_tuser;

  wire [63:0] tx_axis_tdata;
  wire [7:0] tx_axis_tkeep;
  wire tx_axis_tvalid;
  wire tx_axis_tready;
  wire tx_axis_tlast;
  wire tx_axis_tuser;

  wire [511:0] rx_512_axis_tdata;
  wire [63:0] rx_512_axis_tkeep;
  wire rx_512_axis_tvalid;
  wire rx_512_axis_tready;
  wire rx_512_axis_tlast;
  wire rx_512_axis_tuser;

  wire [511:0] tx_512_axis_tdata;
  wire [63:0] tx_512_axis_tkeep;
  wire tx_512_axis_tvalid;
  wire tx_512_axis_tready;
  wire tx_512_axis_tlast;
  wire tx_512_axis_tuser;

  wire [511:0] tx_512_fifo_axis_tdata;
  wire [63:0] tx_512_fifo_axis_tkeep;
  wire tx_512_fifo_axis_tvalid;
  wire tx_512_fifo_axis_tready;
  wire tx_512_fifo_axis_tlast;
  wire tx_512_fifo_axis_tuser;

  // Ethernet frame between Ethernet modules and UDP stack
  wire rx_eth_hdr_ready;
  wire rx_eth_hdr_valid;
  wire [47:0] rx_eth_dest_mac;
  wire [47:0] rx_eth_src_mac;
  wire [15:0] rx_eth_type;
  wire [511:0] rx_eth_payload_axis_tdata;
  wire [63:0] rx_eth_payload_axis_tkeep;
  wire rx_eth_payload_axis_tvalid;
  wire rx_eth_payload_axis_tready;
  wire rx_eth_payload_axis_tlast;
  wire rx_eth_payload_axis_tuser;

  wire tx_eth_hdr_ready;
  wire tx_eth_hdr_valid;
  wire [47:0] tx_eth_dest_mac;
  wire [47:0] tx_eth_src_mac;
  wire [15:0] tx_eth_type;
  wire [511:0] tx_eth_payload_axis_tdata;
  wire [63:0] tx_eth_payload_axis_tkeep;
  wire tx_eth_payload_axis_tvalid;
  wire tx_eth_payload_axis_tready;
  wire tx_eth_payload_axis_tlast;
  wire tx_eth_payload_axis_tuser;

  // IP frame connections
  wire rx_ip_hdr_valid;
  wire rx_ip_hdr_ready;
  wire [47:0] rx_ip_eth_dest_mac;
  wire [47:0] rx_ip_eth_src_mac;
  wire [15:0] rx_ip_eth_type;
  wire [3:0] rx_ip_version;
  wire [3:0] rx_ip_ihl;
  wire [5:0] rx_ip_dscp;
  wire [1:0] rx_ip_ecn;
  wire [15:0] rx_ip_length;
  wire [15:0] rx_ip_identification;
  wire [2:0] rx_ip_flags;
  wire [12:0] rx_ip_fragment_offset;
  wire [7:0] rx_ip_ttl;
  wire [7:0] rx_ip_protocol;
  wire [15:0] rx_ip_header_checksum;
  wire [31:0] rx_ip_source_ip;
  wire [31:0] rx_ip_dest_ip;
  wire [511:0] rx_ip_payload_axis_tdata;
  wire [63:0] rx_ip_payload_axis_tkeep;
  wire rx_ip_payload_axis_tvalid;
  wire rx_ip_payload_axis_tready;
  wire rx_ip_payload_axis_tlast;
  wire rx_ip_payload_axis_tuser;

  wire tx_ip_hdr_valid;
  wire tx_ip_hdr_ready;
  wire [5:0] tx_ip_dscp;
  wire [1:0] tx_ip_ecn;
  wire [15:0] tx_ip_length;
  wire [7:0] tx_ip_ttl;
  wire [7:0] tx_ip_protocol;
  wire [31:0] tx_ip_source_ip;
  wire [31:0] tx_ip_dest_ip;
  wire [511:0] tx_ip_payload_axis_tdata;
  wire [63:0] tx_ip_payload_axis_tkeep;
  wire tx_ip_payload_axis_tvalid;
  wire tx_ip_payload_axis_tready;
  wire tx_ip_payload_axis_tlast;
  wire tx_ip_payload_axis_tuser;

  // UDP frame connections
  wire rx_udp_hdr_valid;
  wire rx_udp_hdr_ready;
  wire [47:0] rx_udp_eth_dest_mac;
  wire [47:0] rx_udp_eth_src_mac;
  wire [15:0] rx_udp_eth_type;
  wire [3:0] rx_udp_ip_version;
  wire [3:0] rx_udp_ip_ihl;
  wire [5:0] rx_udp_ip_dscp;
  wire [1:0] rx_udp_ip_ecn;
  wire [15:0] rx_udp_ip_length;
  wire [15:0] rx_udp_ip_identification;
  wire [2:0] rx_udp_ip_flags;
  wire [12:0] rx_udp_ip_fragment_offset;
  wire [7:0] rx_udp_ip_ttl;
  wire [7:0] rx_udp_ip_protocol;
  wire [15:0] rx_udp_ip_header_checksum;
  wire [31:0] rx_udp_ip_source_ip;
  wire [31:0] rx_udp_ip_dest_ip;
  wire [15:0] rx_udp_source_port;
  wire [15:0] rx_udp_dest_port;
  wire [15:0] rx_udp_length;
  wire [15:0] rx_udp_checksum;
  wire [511:0] rx_udp_payload_axis_tdata;
  wire [63:0] rx_udp_payload_axis_tkeep;
  wire rx_udp_payload_axis_tvalid;
  wire rx_udp_payload_axis_tready;
  wire rx_udp_payload_axis_tlast;
  wire rx_udp_payload_axis_tuser;

  wire tx_udp_hdr_valid;
  wire tx_udp_hdr_ready;
  wire [5:0] tx_udp_ip_dscp;
  wire [1:0] tx_udp_ip_ecn;
  wire [7:0] tx_udp_ip_ttl;
  wire [31:0] tx_udp_ip_source_ip;
  wire [31:0] tx_udp_ip_dest_ip;
  wire [15:0] tx_udp_source_port;
  wire [15:0] tx_udp_dest_port;
  wire [15:0] tx_udp_length;
  wire [15:0] tx_udp_checksum;
  wire [511:0] tx_udp_payload_axis_tdata;
  wire [63:0] tx_udp_payload_axis_tkeep;
  wire tx_udp_payload_axis_tvalid;
  wire tx_udp_payload_axis_tready;
  wire tx_udp_payload_axis_tlast;
  wire tx_udp_payload_axis_tuser;

  wire [511:0] rx_fifo_udp_payload_axis_tdata;
  wire [63:0] rx_fifo_udp_payload_axis_tkeep;
  wire rx_fifo_udp_payload_axis_tvalid;
  wire rx_fifo_udp_payload_axis_tready;
  wire rx_fifo_udp_payload_axis_tlast;
  wire rx_fifo_udp_payload_axis_tuser;

  wire [511:0] tx_fifo_udp_payload_axis_tdata;
  wire [63:0] tx_fifo_udp_payload_axis_tkeep;
  wire tx_fifo_udp_payload_axis_tvalid;
  wire tx_fifo_udp_payload_axis_tready;
  wire tx_fifo_udp_payload_axis_tlast;
  wire tx_fifo_udp_payload_axis_tuser;

  // Configuration
  wire [47:0] local_mac   = 48'h02_00_00_00_00_00;
  wire [31:0] local_ip    = {8'd22 , 8'd1  , 8'd212, 8'd10};
  wire [31:0] dest_ip     = {8'd22 , 8'd1  , 8'd212, 8'd11};
  wire [31:0] gateway_ip  = {8'd22 , 8'd1  , 8'd212,  8'd1};
  wire [31:0] subnet_mask = {8'd255, 8'd255, 8'd255,  8'd0};

  // IP ports not used
  assign rx_ip_hdr_ready = 1;
  assign rx_ip_payload_axis_tready = 1;

  assign tx_ip_hdr_valid = 0;
  assign tx_ip_dscp = 0;
  assign tx_ip_ecn = 0;
  assign tx_ip_length = 0;
  assign tx_ip_ttl = 0;
  assign tx_ip_protocol = 0;
  assign tx_ip_source_ip = 0;
  assign tx_ip_dest_ip = 0;
  assign tx_ip_payload_axis_tdata = 0;
  assign tx_ip_payload_axis_tkeep = 0;
  assign tx_ip_payload_axis_tvalid = 0;
  assign tx_ip_payload_axis_tlast = 0;
  assign tx_ip_payload_axis_tuser = 0;

  // Loop back UDP
  wire match_cond = rx_udp_dest_port == 1234;
  wire no_match = !match_cond;

  reg match_cond_reg = 0;
  reg no_match_reg = 0;

  always @(posedge clk) begin
    if (rst) begin
      match_cond_reg <= 0;
      no_match_reg   <= 0;
    end else begin
      if (rx_udp_payload_axis_tvalid) begin
        if ((!match_cond_reg && !no_match_reg) ||
                (rx_udp_payload_axis_tvalid && rx_udp_payload_axis_tready && rx_udp_payload_axis_tlast)) begin
          match_cond_reg <= match_cond;
          no_match_reg   <= no_match;
        end
      end else begin
        match_cond_reg <= 0;
        no_match_reg   <= 0;
      end
    end
  end

  /*
  assign tx_udp_hdr_valid = rx_udp_hdr_valid && match_cond;
  assign rx_udp_hdr_ready = (tx_eth_hdr_ready && match_cond) || no_match;
  assign tx_udp_ip_dscp = 0;
  assign tx_udp_ip_ecn = 0;
  assign tx_udp_ip_ttl = 64;
  assign tx_udp_ip_source_ip = local_ip;
  assign tx_udp_ip_dest_ip = rx_udp_ip_source_ip;
  assign tx_udp_source_port = rx_udp_dest_port;
  assign tx_udp_dest_port = rx_udp_source_port;
  assign tx_udp_length = rx_udp_length;
  assign tx_udp_checksum = 0;

  assign tx_udp_payload_axis_tdata = tx_fifo_udp_payload_axis_tdata;
  assign tx_udp_payload_axis_tkeep = tx_fifo_udp_payload_axis_tkeep;
  assign tx_udp_payload_axis_tvalid = tx_fifo_udp_payload_axis_tvalid;
  assign tx_fifo_udp_payload_axis_tready = tx_udp_payload_axis_tready;
  assign tx_udp_payload_axis_tlast = tx_fifo_udp_payload_axis_tlast;
  assign tx_udp_payload_axis_tuser = tx_fifo_udp_payload_axis_tuser;
  */
  /*
  assign rx_fifo_udp_payload_axis_tdata = rx_udp_payload_axis_tdata;
  assign rx_fifo_udp_payload_axis_tkeep = rx_udp_payload_axis_tkeep;
  assign rx_fifo_udp_payload_axis_tvalid = rx_udp_payload_axis_tvalid && match_cond_reg;
  assign rx_udp_payload_axis_tready = (rx_fifo_udp_payload_axis_tready && match_cond_reg) || no_match_reg;
  assign rx_fifo_udp_payload_axis_tlast = rx_udp_payload_axis_tlast;
  assign rx_fifo_udp_payload_axis_tuser = rx_udp_payload_axis_tuser;

  */
  // Place first payload byte onto LEDs
  reg valid_last = 0;
  reg [7:0] led_reg = 0;

  always @(posedge clk) begin
    if (rst) begin
      led_reg <= 0;
    end else begin
      valid_last <= tx_udp_payload_axis_tvalid;
      if (tx_udp_payload_axis_tvalid && !valid_last) begin
        led_reg <= tx_udp_payload_axis_tdata;
      end
    end
  end

  //assign led = sw;
  assign led = led_reg;
  //assign phy_reset_n = !rst;

  eth_mac_10g_fifo #(
      .ENABLE_PADDING(1),
      .ENABLE_DIC(1),
      .MIN_FRAME_LENGTH(64),
      .TX_FIFO_DEPTH(4096),
      .TX_FRAME_FIFO(1),
      .RX_FIFO_DEPTH(4096),
      .RX_FRAME_FIFO(1)
  ) eth_mac_10g_fifo_inst (
      .rx_clk(xgmii_rx_clk),
      .rx_rst(xgmii_rx_rst),
      .tx_clk(xgmii_tx_clk),
      .tx_rst(xgmii_tx_rst),
      .logic_clk(clk),
      .logic_rst(rst),

      .tx_axis_tdata (tx_axis_tdata),
      .tx_axis_tkeep (tx_axis_tkeep),
      .tx_axis_tvalid(tx_axis_tvalid),
      .tx_axis_tready(tx_axis_tready),
      .tx_axis_tlast (tx_axis_tlast),
      .tx_axis_tuser (tx_axis_tuser),

      .rx_axis_tdata (rx_axis_tdata),
      .rx_axis_tkeep (rx_axis_tkeep),
      .rx_axis_tvalid(rx_axis_tvalid),
      .rx_axis_tready(rx_axis_tready),
      .rx_axis_tlast (rx_axis_tlast),
      .rx_axis_tuser (rx_axis_tuser),

      .xgmii_rxd(xgmii_rxd),
      .xgmii_rxc(xgmii_rxc),
      .xgmii_txd(xgmii_txd),
      .xgmii_txc(xgmii_txc),

      .tx_fifo_overflow  (),
      .tx_fifo_bad_frame (),
      .tx_fifo_good_frame(),
      .rx_error_bad_frame(),
      .rx_error_bad_fcs  (),
      .rx_fifo_overflow  (),
      .rx_fifo_bad_frame (),
      .rx_fifo_good_frame(),

      .cfg_ifg(8'd12),
      .cfg_tx_enable(1'b1),
      .cfg_rx_enable(1'b1)
  );


  // tap port mux logic
  // sw[3] enable
  // sw[2] select 0 rx, 1 tx

  reg [1:0] mac_rx_tdest;
  reg [1:0] tx_tdest;
  reg [1:0] gig_rx_tdest;

  always @* begin
    if (sw[3]) begin
      if (sw[2]) begin
        // Tap on TX path
        // MAC RX out -> stack RX in
        // stack TX out -> gig TX in
        // gig RX out -> MAC TX in
        mac_rx_tdest = 2'd1;
        tx_tdest = 2'd2;
        gig_rx_tdest = 2'd0;
      end else begin
        // Tap on RX path
        // MAC RX out -> gig TX in
        // stack TX out -> MAC TX in
        // gig RX out -> stack RX in
        mac_rx_tdest = 2'd2;
        tx_tdest = 2'd0;
        gig_rx_tdest = 2'd1;
      end
    end else begin
      // Tap disabled
      // MAC RX out -> stack RX in
      // stack TX out -> MAC TX in
      // gig RX out -> blackhole
      mac_rx_tdest = 2'd1;
      tx_tdest = 2'd0;
      gig_rx_tdest = 2'd3;
    end
  end

  axis_adapter #(
      .S_DATA_WIDTH(64),
      .M_DATA_WIDTH(512),
      .ID_ENABLE(0),
      .DEST_ENABLE(0),
      .USER_ENABLE(1),
      .USER_WIDTH(1)
  ) rx_axis_64_to_512_adapter_inst (
      .clk(clk),
      .rst(rst),
      // AXI input
      .s_axis_tdata(rx_axis_tdata),
      .s_axis_tkeep(rx_axis_tkeep),
      .s_axis_tvalid(rx_axis_tvalid),
      .s_axis_tready(rx_axis_tready),
      .s_axis_tlast(rx_axis_tlast),
      .s_axis_tuser(rx_axis_tuser),
      // AXI output
      .m_axis_tdata(rx_512_axis_tdata),
      .m_axis_tkeep(rx_512_axis_tkeep),
      .m_axis_tvalid(rx_512_axis_tvalid),
      .m_axis_tready(rx_512_axis_tready),
      .m_axis_tlast(rx_512_axis_tlast),
      .m_axis_tuser(rx_512_axis_tuser)
  );

  axis_adapter #(
      .S_DATA_WIDTH(512),
      .M_DATA_WIDTH(64),
      .ID_ENABLE(0),
      .DEST_ENABLE(0),
      .USER_ENABLE(1),
      .USER_WIDTH(1)
  ) tx_axis_512_to_64_adapter_inst (
      .clk(clk),
      .rst(rst),
      // AXI input
      .s_axis_tdata(tx_512_axis_tdata),
      .s_axis_tkeep(tx_512_axis_tkeep),
      .s_axis_tvalid(tx_512_axis_tvalid),
      .s_axis_tready(tx_512_axis_tready),
      .s_axis_tlast(tx_512_axis_tlast),
      .s_axis_tuser(tx_512_axis_tuser),
      // AXI output
      .m_axis_tdata(tx_axis_tdata),
      .m_axis_tkeep(tx_axis_tkeep),
      .m_axis_tvalid(tx_axis_tvalid),
      .m_axis_tready(tx_axis_tready),
      .m_axis_tlast(tx_axis_tlast),
      .m_axis_tuser(tx_axis_tuser)
  );


  eth_axis_rx #(
      .DATA_WIDTH(512)
  ) eth_axis_rx_inst (
      .clk(clk),
      .rst(rst),
      // AXI input
      .s_axis_tdata(rx_512_axis_tdata),
      .s_axis_tkeep(rx_512_axis_tkeep),
      .s_axis_tvalid(rx_512_axis_tvalid),
      .s_axis_tready(rx_512_axis_tready),
      .s_axis_tlast(rx_512_axis_tlast),
      .s_axis_tuser(rx_512_axis_tuser),
      // Ethernet frame output
      .m_eth_hdr_valid(rx_eth_hdr_valid),
      .m_eth_hdr_ready(rx_eth_hdr_ready),
      .m_eth_dest_mac(rx_eth_dest_mac),
      .m_eth_src_mac(rx_eth_src_mac),
      .m_eth_type(rx_eth_type),
      .m_eth_payload_axis_tdata(rx_eth_payload_axis_tdata),
      .m_eth_payload_axis_tkeep(rx_eth_payload_axis_tkeep),
      .m_eth_payload_axis_tvalid(rx_eth_payload_axis_tvalid),
      .m_eth_payload_axis_tready(rx_eth_payload_axis_tready),
      .m_eth_payload_axis_tlast(rx_eth_payload_axis_tlast),
      .m_eth_payload_axis_tuser(rx_eth_payload_axis_tuser),
      // Status signals
      .busy(),
      .error_header_early_termination()
  );

  eth_axis_tx #(
      .DATA_WIDTH(512)
  ) eth_axis_tx_inst (
      .clk                      (clk),
      .rst                      (rst),
      // Ethernet frame input
      .s_eth_hdr_valid          (tx_eth_hdr_valid),
      .s_eth_hdr_ready          (tx_eth_hdr_ready),
      .s_eth_dest_mac           (tx_eth_dest_mac),
      .s_eth_src_mac            (tx_eth_src_mac),
      .s_eth_type               (tx_eth_type),
      .s_eth_payload_axis_tdata (tx_eth_payload_axis_tdata),
      .s_eth_payload_axis_tkeep (tx_eth_payload_axis_tkeep),
      .s_eth_payload_axis_tvalid(tx_eth_payload_axis_tvalid),
      .s_eth_payload_axis_tready(tx_eth_payload_axis_tready),
      .s_eth_payload_axis_tlast (tx_eth_payload_axis_tlast),
      .s_eth_payload_axis_tuser (tx_eth_payload_axis_tuser),
      // AXI output
      .m_axis_tdata             (tx_512_fifo_axis_tdata),
      .m_axis_tkeep             (tx_512_fifo_axis_tkeep),
      .m_axis_tvalid            (tx_512_fifo_axis_tvalid),
      .m_axis_tready            (tx_512_fifo_axis_tready),
      .m_axis_tlast             (tx_512_fifo_axis_tlast),
      .m_axis_tuser             (tx_512_fifo_axis_tuser),
      // Status signals
      .busy                     ()
  );

  axis_fifo #(
      .DEPTH(2048),
      .DATA_WIDTH(512),
      .KEEP_ENABLE(1),
      .KEEP_WIDTH(64),
      .ID_ENABLE(0),
      .DEST_ENABLE(0),
      .USER_ENABLE(1),
      .USER_WIDTH(1),
      .FRAME_FIFO(0)
  ) eth_tx_axis_fifo (
      .clk(clk),
      .rst(rst),

      // AXI input
      .s_axis_tdata(tx_512_fifo_axis_tdata),
      .s_axis_tkeep(tx_512_fifo_axis_tkeep),
      .s_axis_tvalid(tx_512_fifo_axis_tvalid),
      .s_axis_tready(tx_512_fifo_axis_tready),
      .s_axis_tlast(tx_512_fifo_axis_tlast),
      .s_axis_tid(0),
      .s_axis_tdest(0),
      .s_axis_tuser(tx_512_fifo_axis_tuser),

      // AXI output
      .m_axis_tdata(tx_512_axis_tdata),
      .m_axis_tkeep(tx_512_axis_tkeep),
      .m_axis_tvalid(tx_512_axis_tvalid),
      .m_axis_tready(tx_512_axis_tready),
      .m_axis_tlast(tx_512_axis_tlast),
      .m_axis_tid(),
      .m_axis_tdest(),
      .m_axis_tuser(tx_512_axis_tuser),

      // Status
      .status_overflow  (),
      .status_bad_frame (),
      .status_good_frame()
  );

  udp_complete_512 #(
      .UDP_CHECKSUM_GEN_ENABLE(0)
  ) udp_complete_inst (
      .clk(clk),
      .rst(rst),
      // Ethernet frame input
      .s_eth_hdr_valid(rx_eth_hdr_valid),
      .s_eth_hdr_ready(rx_eth_hdr_ready),
      .s_eth_dest_mac(rx_eth_dest_mac),
      .s_eth_src_mac(rx_eth_src_mac),
      .s_eth_type(rx_eth_type),
      .s_eth_payload_axis_tdata(rx_eth_payload_axis_tdata),
      .s_eth_payload_axis_tkeep(rx_eth_payload_axis_tkeep),
      .s_eth_payload_axis_tvalid(rx_eth_payload_axis_tvalid),
      .s_eth_payload_axis_tready(rx_eth_payload_axis_tready),
      .s_eth_payload_axis_tlast(rx_eth_payload_axis_tlast),
      .s_eth_payload_axis_tuser(rx_eth_payload_axis_tuser),
      // Ethernet frame output
      .m_eth_hdr_valid(tx_eth_hdr_valid),
      .m_eth_hdr_ready(tx_eth_hdr_ready),
      .m_eth_dest_mac(tx_eth_dest_mac),
      .m_eth_src_mac(tx_eth_src_mac),
      .m_eth_type(tx_eth_type),
      .m_eth_payload_axis_tdata(tx_eth_payload_axis_tdata),
      .m_eth_payload_axis_tkeep(tx_eth_payload_axis_tkeep),
      .m_eth_payload_axis_tvalid(tx_eth_payload_axis_tvalid),
      .m_eth_payload_axis_tready(tx_eth_payload_axis_tready),
      .m_eth_payload_axis_tlast(tx_eth_payload_axis_tlast),
      .m_eth_payload_axis_tuser(tx_eth_payload_axis_tuser),
      // IP frame input
      .s_ip_hdr_valid(tx_ip_hdr_valid),
      .s_ip_hdr_ready(tx_ip_hdr_ready),
      .s_ip_dscp(tx_ip_dscp),
      .s_ip_ecn(tx_ip_ecn),
      .s_ip_length(tx_ip_length),
      .s_ip_ttl(tx_ip_ttl),
      .s_ip_protocol(tx_ip_protocol),
      .s_ip_source_ip(tx_ip_source_ip),
      .s_ip_dest_ip(tx_ip_dest_ip),
      .s_ip_payload_axis_tdata(tx_ip_payload_axis_tdata),
      .s_ip_payload_axis_tkeep(tx_ip_payload_axis_tkeep),
      .s_ip_payload_axis_tvalid(tx_ip_payload_axis_tvalid),
      .s_ip_payload_axis_tready(tx_ip_payload_axis_tready),
      .s_ip_payload_axis_tlast(tx_ip_payload_axis_tlast),
      .s_ip_payload_axis_tuser(tx_ip_payload_axis_tuser),
      // IP frame output
      .m_ip_hdr_valid(rx_ip_hdr_valid),
      .m_ip_hdr_ready(rx_ip_hdr_ready),
      .m_ip_eth_dest_mac(rx_ip_eth_dest_mac),
      .m_ip_eth_src_mac(rx_ip_eth_src_mac),
      .m_ip_eth_type(rx_ip_eth_type),
      .m_ip_version(rx_ip_version),
      .m_ip_ihl(rx_ip_ihl),
      .m_ip_dscp(rx_ip_dscp),
      .m_ip_ecn(rx_ip_ecn),
      .m_ip_length(rx_ip_length),
      .m_ip_identification(rx_ip_identification),
      .m_ip_flags(rx_ip_flags),
      .m_ip_fragment_offset(rx_ip_fragment_offset),
      .m_ip_ttl(rx_ip_ttl),
      .m_ip_protocol(rx_ip_protocol),
      .m_ip_header_checksum(rx_ip_header_checksum),
      .m_ip_source_ip(rx_ip_source_ip),
      .m_ip_dest_ip(rx_ip_dest_ip),
      .m_ip_payload_axis_tdata(rx_ip_payload_axis_tdata),
      .m_ip_payload_axis_tkeep(rx_ip_payload_axis_tkeep),
      .m_ip_payload_axis_tvalid(rx_ip_payload_axis_tvalid),
      .m_ip_payload_axis_tready(rx_ip_payload_axis_tready),
      .m_ip_payload_axis_tlast(rx_ip_payload_axis_tlast),
      .m_ip_payload_axis_tuser(rx_ip_payload_axis_tuser),
      // UDP frame input
      .s_udp_hdr_valid(tx_udp_hdr_valid),
      .s_udp_hdr_ready(tx_udp_hdr_ready),
      .s_udp_ip_dscp(tx_udp_ip_dscp),
      .s_udp_ip_ecn(tx_udp_ip_ecn),
      .s_udp_ip_ttl(tx_udp_ip_ttl),
      .s_udp_ip_source_ip(tx_udp_ip_source_ip),
      .s_udp_ip_dest_ip(tx_udp_ip_dest_ip),
      .s_udp_source_port(tx_udp_source_port),
      .s_udp_dest_port(tx_udp_dest_port),
      .s_udp_length(tx_udp_length),
      .s_udp_checksum(tx_udp_checksum),
      .s_udp_payload_axis_tdata(tx_udp_payload_axis_tdata),
      .s_udp_payload_axis_tkeep(tx_udp_payload_axis_tkeep),
      .s_udp_payload_axis_tvalid(tx_udp_payload_axis_tvalid),
      .s_udp_payload_axis_tready(tx_udp_payload_axis_tready),
      .s_udp_payload_axis_tlast(tx_udp_payload_axis_tlast),
      .s_udp_payload_axis_tuser(tx_udp_payload_axis_tuser),
      // UDP frame output
      .m_udp_hdr_valid(rx_udp_hdr_valid),
      .m_udp_hdr_ready(rx_udp_hdr_ready),
      .m_udp_eth_dest_mac(rx_udp_eth_dest_mac),
      .m_udp_eth_src_mac(rx_udp_eth_src_mac),
      .m_udp_eth_type(rx_udp_eth_type),
      .m_udp_ip_version(rx_udp_ip_version),
      .m_udp_ip_ihl(rx_udp_ip_ihl),
      .m_udp_ip_dscp(rx_udp_ip_dscp),
      .m_udp_ip_ecn(rx_udp_ip_ecn),
      .m_udp_ip_length(rx_udp_ip_length),
      .m_udp_ip_identification(rx_udp_ip_identification),
      .m_udp_ip_flags(rx_udp_ip_flags),
      .m_udp_ip_fragment_offset(rx_udp_ip_fragment_offset),
      .m_udp_ip_ttl(rx_udp_ip_ttl),
      .m_udp_ip_protocol(rx_udp_ip_protocol),
      .m_udp_ip_header_checksum(rx_udp_ip_header_checksum),
      .m_udp_ip_source_ip(rx_udp_ip_source_ip),
      .m_udp_ip_dest_ip(rx_udp_ip_dest_ip),
      .m_udp_source_port(rx_udp_source_port),
      .m_udp_dest_port(rx_udp_dest_port),
      .m_udp_length(rx_udp_length),
      .m_udp_checksum(rx_udp_checksum),
      .m_udp_payload_axis_tdata(rx_udp_payload_axis_tdata),
      .m_udp_payload_axis_tkeep(rx_udp_payload_axis_tkeep),
      .m_udp_payload_axis_tvalid(rx_udp_payload_axis_tvalid),
      .m_udp_payload_axis_tready(rx_udp_payload_axis_tready),
      .m_udp_payload_axis_tlast(rx_udp_payload_axis_tlast),
      .m_udp_payload_axis_tuser(rx_udp_payload_axis_tuser),
      // Status signals
      .ip_rx_busy(),
      .ip_tx_busy(),
      .udp_rx_busy(),
      .udp_tx_busy(),
      .ip_rx_error_header_early_termination(),
      .ip_rx_error_payload_early_termination(),
      .ip_rx_error_invalid_header(),
      .ip_rx_error_invalid_checksum(),
      .ip_tx_error_payload_early_termination(),
      .ip_tx_error_arp_failed(),
      .udp_rx_error_header_early_termination(),
      .udp_rx_error_payload_early_termination(),
      .udp_tx_error_payload_early_termination(),
      // Configuration
      .local_mac(local_mac),
      .local_ip(local_ip),
      .gateway_ip(gateway_ip),
      .subnet_mask(subnet_mask),
      .clear_arp_cache(1'b0)
  );

  assign rx_fifo_udp_payload_axis_tready = 1'b1;


  wire [31:0] dma_transfer_length;
  wire [23:0] rem_qpn;
  wire [23:0] rem_psn;
  wire [31:0] r_key;
  wire [47:0] rem_addr;
  wire [31:0] rem_ip_addr = {8'd22, 8'd1, 8'd212, 8'd11};
  wire start_transfer;

  wire metadata_valid;

  // ROCE TX inst
  RoCE_minimal_stack_512 RoCE_minimal_stack_512_instance (
      .clk(clk),
      .rst(rst),
      .s_udp_hdr_valid(rx_udp_hdr_valid),
      .s_udp_hdr_ready(rx_udp_hdr_ready),
      .s_eth_dest_mac(rx_udp_eth_dest_mac),
      .s_eth_src_mac(rx_udp_eth_src_mac),
      .s_eth_type(rx_udp_eth_type),
      .s_ip_version(rx_udp_ip_version),
      .s_ip_ihl(rx_udp_ip_ihl),
      .s_ip_dscp(rx_udp_ip_dscp),
      .s_ip_ecn(rx_udp_ip_ecn),
      .s_ip_length(rx_udp_ip_length),
      .s_ip_identification(rx_udp_ip_identification),
      .s_ip_flags(rx_udp_ip_flags),
      .s_ip_fragment_offset(rx_udp_ip_fragment_offset),
      .s_ip_ttl(rx_udp_ip_ttl),
      .s_ip_protocol(rx_udp_ip_protocol),
      .s_ip_header_checksum(rx_udp_ip_header_checksum),
      .s_ip_source_ip(rx_udp_ip_source_ip),
      .s_ip_dest_ip(rx_udp_ip_dest_ip),
      .s_udp_source_port(rx_udp_source_port),
      .s_udp_dest_port(rx_udp_dest_port),
      .s_udp_length(rx_udp_length),
      .s_udp_checksum(rx_udp_checksum),
      .s_udp_payload_axis_tdata(rx_udp_payload_axis_tdata),
      .s_udp_payload_axis_tkeep(rx_udp_payload_axis_tkeep),
      .s_udp_payload_axis_tvalid(rx_udp_payload_axis_tvalid),
      .s_udp_payload_axis_tready(rx_udp_payload_axis_tready),
      .s_udp_payload_axis_tlast(rx_udp_payload_axis_tlast),
      .s_udp_payload_axis_tuser(rx_udp_payload_axis_tuser),
      .m_udp_hdr_valid(tx_udp_hdr_valid),
      .m_udp_hdr_ready(tx_udp_hdr_ready),
      .m_eth_dest_mac(),
      .m_eth_src_mac(),
      .m_eth_type(),
      .m_ip_version(),
      .m_ip_ihl(),
      .m_ip_dscp(tx_udp_ip_dscp),
      .m_ip_ecn(tx_udp_ip_ecn),
      .m_ip_length(),
      .m_ip_identification(),
      .m_ip_flags(),
      .m_ip_fragment_offset(),
      .m_ip_ttl(tx_udp_ip_ttl),
      .m_ip_protocol(),
      .m_ip_header_checksum(),
      .m_ip_source_ip(tx_udp_ip_source_ip),
      .m_ip_dest_ip(tx_udp_ip_dest_ip),
      .m_udp_source_port(tx_udp_source_port),
      .m_udp_dest_port(tx_udp_dest_port),
      .m_udp_length(tx_udp_length),
      .m_udp_checksum(tx_udp_checksum),
      .m_udp_payload_axis_tdata(tx_udp_payload_axis_tdata),
      .m_udp_payload_axis_tkeep(tx_udp_payload_axis_tkeep),
      .m_udp_payload_axis_tvalid(tx_udp_payload_axis_tvalid),
      .m_udp_payload_axis_tready(tx_udp_payload_axis_tready),
      .m_udp_payload_axis_tlast(tx_udp_payload_axis_tlast),
      .m_udp_payload_axis_tuser(tx_udp_payload_axis_tuser),
      .busy(),
      .error_payload_early_termination(),
      .pmtu(13'd2048),
      .RoCE_udp_port(16'h12B7),
      .loc_ip_addr(local_ip)
  );

  /*
axis_fifo #(
    .DEPTH(8192),
    .DATA_WIDTH(64),
    .KEEP_ENABLE(1),
    .KEEP_WIDTH(8),
    .ID_ENABLE(0),
    .DEST_ENABLE(0),
    .USER_ENABLE(1),
    .USER_WIDTH(1),
    .FRAME_FIFO(0)
)
udp_payload_fifo (
    .clk(clk),
    .rst(rst),

    // AXI input
    .s_axis_tdata(rx_fifo_udp_payload_axis_tdata),
    .s_axis_tkeep(rx_fifo_udp_payload_axis_tkeep),
    .s_axis_tvalid(rx_fifo_udp_payload_axis_tvalid),
    .s_axis_tready(rx_fifo_udp_payload_axis_tready),
    .s_axis_tlast(rx_fifo_udp_payload_axis_tlast),
    .s_axis_tid(0),
    .s_axis_tdest(0),
    .s_axis_tuser(rx_fifo_udp_payload_axis_tuser),

    // AXI output
    .m_axis_tdata(tx_fifo_udp_payload_axis_tdata),
    .m_axis_tkeep(tx_fifo_udp_payload_axis_tkeep),
    .m_axis_tvalid(tx_fifo_udp_payload_axis_tvalid),
    .m_axis_tready(tx_fifo_udp_payload_axis_tready),
    .m_axis_tlast(tx_fifo_udp_payload_axis_tlast),
    .m_axis_tid(),
    .m_axis_tdest(),
    .m_axis_tuser(tx_fifo_udp_payload_axis_tuser),

    // Status
    .status_overflow(),
    .status_bad_frame(),
    .status_good_frame()
);

*/
endmodule

`resetall
