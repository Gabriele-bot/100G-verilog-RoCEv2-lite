`timescale 1ns / 1ps

package Board_params;

    parameter RoCE_CLOCK_PERIOD = 1000/156.25; // in ns
    parameter MAC_CLOCK_PERIOD = 1000/156.25; // in ns
  
endpackage
