package Board_params;

    parameter NET_CLOCK_PERIOD = 6.4; // in ns
    parameter MAC_CLOCK_PERIOD = 6.4; // in ns

    parameter NET_DATA_WIDTH = 512;
  
endpackage
