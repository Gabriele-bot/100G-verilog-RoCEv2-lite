library IEEE;
use IEEE.std_logic_1164.all;

entity CRC32_D512_pipeline_with_keep is
    generic(
        REVERSE_INPUT  : boolean                       := FALSE;
        REVERSE_RESULT : boolean                       := FALSE;
        FINXOR         : std_logic_vector(31 downto 0) := X"00000000"
    );
    port(
        clk           : in  std_logic;
        rst           : in  std_logic;
        crcIn         : in  std_logic_vector(31 downto 0);
        data_in       : in  std_logic_vector(511 downto 0);
        keep_in       : in  std_logic_vector(63 downto 0);
        valid_in      : in  std_logic;
        crcOut        : out std_logic_vector(31 downto 0);
        valid_crc_out : out std_logic
    );
end entity CRC32_D512_pipeline_with_keep;

architecture Behavioral of CRC32_D512_pipeline_with_keep is

    type crc_pipeline_stage_t is array (15 downto 0) of std_logic_vector(31 downto 0);
    signal crc_stage : crc_pipeline_stage_t;

    type data_pipeline_stage_t is array (16 downto 0) of std_logic_vector(511 downto 0);
    signal data_stage : data_pipeline_stage_t;

    type keep_pipeline_stage_t is array (16 downto 0) of std_logic_vector(63 downto 0);
    signal keep_stage : keep_pipeline_stage_t;

    signal valid_shreg : std_logic_vector(16 downto 0);

    signal data : std_logic_vector(511 downto 0);

    signal crc_rev : std_logic_vector(31 downto 0);

begin

    reverse_in_g : if REVERSE_INPUT generate
        reverse_g : for i in 0 to 511 generate
            data(i) <= data_in(511 - i);
        end generate;
    else generate
        data <= data_in;
    end generate;

    valid_shreg(0) <= valid_in;
    process(clk)
    begin
        if rising_edge(clk) then
            valid_shreg(valid_shreg'high downto 1) <= valid_shreg(valid_shreg'high - 1 downto 0);
        end if;
    end process;

    data_stage(0) <= data;
    process(clk)
    begin
        if rising_edge(clk) then
            data_stage(data_stage'high downto 1) <= data_stage(data_stage'high - 1 downto 0);
        end if;
    end process;

    keep_stage(0) <= keep_in;
    process(clk)
    begin
        if rising_edge(clk) then
            keep_stage(keep_stage'high downto 1) <= keep_stage(keep_stage'high - 1 downto 0);
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(0)(3 downto 0) = X"F" then
                crc_stage(0)(0)  <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(12) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(26) xor data_stage(0)(29) xor data_stage(0)(30) xor data_stage(0)(31);
                crc_stage(0)(1)  <= data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(7) xor data_stage(0)(11) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(27) xor data_stage(0)(30) xor data_stage(0)(31);
                crc_stage(0)(2)  <= data_stage(0)(0) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(6) xor data_stage(0)(7) xor data_stage(0)(8) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(28) xor data_stage(0)(31);
                crc_stage(0)(3)  <= data_stage(0)(1) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(7) xor data_stage(0)(8) xor data_stage(0)(9) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(27) xor data_stage(0)(29);
                crc_stage(0)(4)  <= data_stage(0)(0) xor data_stage(0)(2) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(27) xor data_stage(0)(28) xor data_stage(0)(30);
                crc_stage(0)(5)  <= data_stage(0)(1) xor data_stage(0)(3) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(27) xor data_stage(0)(28) xor data_stage(0)(29) xor data_stage(0)(31);
                crc_stage(0)(6)  <= data_stage(0)(1) xor data_stage(0)(5) xor data_stage(0)(7) xor data_stage(0)(8) xor data_stage(0)(16) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(25) xor data_stage(0)(27) xor data_stage(0)(28) xor data_stage(0)(31);
                crc_stage(0)(7)  <= data_stage(0)(0) xor data_stage(0)(2) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(9) xor data_stage(0)(17) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(26) xor data_stage(0)(28) xor data_stage(0)(29);
                crc_stage(0)(8)  <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(3) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(18) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(27) xor data_stage(0)(29) xor data_stage(0)(30);
                crc_stage(0)(9)  <= data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(12) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(28) xor data_stage(0)(29);
                crc_stage(0)(10) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(17) xor data_stage(0)(20) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(27) xor data_stage(0)(31);
                crc_stage(0)(11) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(18) xor data_stage(0)(21) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(28);
                crc_stage(0)(12) <= data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(6) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(11) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(19) xor data_stage(0)(22) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(29);
                crc_stage(0)(13) <= data_stage(0)(0) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(7) xor data_stage(0)(8) xor data_stage(0)(10) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(20) xor data_stage(0)(23) xor data_stage(0)(26) xor data_stage(0)(27) xor data_stage(0)(30);
                crc_stage(0)(14) <= data_stage(0)(1) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(9) xor data_stage(0)(11) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(21) xor data_stage(0)(24) xor data_stage(0)(27) xor data_stage(0)(28) xor data_stage(0)(31);
                crc_stage(0)(15) <= data_stage(0)(2) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(12) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(22) xor data_stage(0)(25) xor data_stage(0)(28) xor data_stage(0)(29);
                crc_stage(0)(16) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(7) xor data_stage(0)(8) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(24) xor data_stage(0)(31);
                crc_stage(0)(17) <= data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(8) xor data_stage(0)(9) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(25);
                crc_stage(0)(18) <= data_stage(0)(0) xor data_stage(0)(2) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(26);
                crc_stage(0)(19) <= data_stage(0)(1) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(7) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(27);
                crc_stage(0)(20) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(7) xor data_stage(0)(8) xor data_stage(0)(10) xor data_stage(0)(16) xor data_stage(0)(18) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(25) xor data_stage(0)(28) xor data_stage(0)(29) xor data_stage(0)(30) xor data_stage(0)(31);
                crc_stage(0)(21) <= data_stage(0)(0) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(12) xor data_stage(0)(18) xor data_stage(0)(20) xor data_stage(0)(21);
                crc_stage(0)(22) <= data_stage(0)(2) xor data_stage(0)(4) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(20) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(26) xor data_stage(0)(29) xor data_stage(0)(30) xor data_stage(0)(31);
                crc_stage(0)(23) <= data_stage(0)(3) xor data_stage(0)(5) xor data_stage(0)(8) xor data_stage(0)(10) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(21) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(27) xor data_stage(0)(30) xor data_stage(0)(31);
                crc_stage(0)(24) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(5) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(12) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(21) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(28) xor data_stage(0)(29) xor data_stage(0)(30);
                crc_stage(0)(25) <= data_stage(0)(0) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(12) xor data_stage(0)(13) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(23) xor data_stage(0)(25);
                crc_stage(0)(26) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(6) xor data_stage(0)(13) xor data_stage(0)(14) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(24) xor data_stage(0)(26);
                crc_stage(0)(27) <= data_stage(0)(0) xor data_stage(0)(4) xor data_stage(0)(7) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(12) xor data_stage(0)(14) xor data_stage(0)(15) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(27) xor data_stage(0)(29) xor data_stage(0)(30) xor data_stage(0)(31);
                crc_stage(0)(28) <= data_stage(0)(2) xor data_stage(0)(4) xor data_stage(0)(6) xor data_stage(0)(8) xor data_stage(0)(10) xor data_stage(0)(13) xor data_stage(0)(15) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(27) xor data_stage(0)(28) xor data_stage(0)(29);
                crc_stage(0)(29) <= data_stage(0)(3) xor data_stage(0)(5) xor data_stage(0)(7) xor data_stage(0)(9) xor data_stage(0)(11) xor data_stage(0)(14) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(26) xor data_stage(0)(28) xor data_stage(0)(29) xor data_stage(0)(30);
                crc_stage(0)(30) <= data_stage(0)(1) xor data_stage(0)(2) xor data_stage(0)(5) xor data_stage(0)(8) xor data_stage(0)(11) xor data_stage(0)(15) xor data_stage(0)(23) xor data_stage(0)(24) xor data_stage(0)(25) xor data_stage(0)(27);
                crc_stage(0)(31) <= data_stage(0)(0) xor data_stage(0)(1) xor data_stage(0)(3) xor data_stage(0)(4) xor data_stage(0)(5) xor data_stage(0)(9) xor data_stage(0)(10) xor data_stage(0)(11) xor data_stage(0)(16) xor data_stage(0)(17) xor data_stage(0)(18) xor data_stage(0)(19) xor data_stage(0)(20) xor data_stage(0)(21) xor data_stage(0)(22) xor data_stage(0)(23) xor data_stage(0)(25) xor data_stage(0)(28) xor data_stage(0)(29) xor data_stage(0)(30) xor data_stage(0)(31);
            else                        --this shuld never happen
                crc_stage(0) <= X"FFFFFFFF";
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(1)(7 downto 4) = X"F" then
                crc_stage(1)(0)  <= crc_stage(0)(0) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(40) xor data_stage(1)(42) xor data_stage(1)(44) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(54) xor data_stage(1)(60) xor data_stage(1)(62) xor data_stage(1)(63);
                crc_stage(1)(1)  <= crc_stage(0)(1) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(41) xor data_stage(1)(43) xor data_stage(1)(45) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(55) xor data_stage(1)(61) xor data_stage(1)(63);
                crc_stage(1)(2)  <= crc_stage(0)(2) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(42) xor data_stage(1)(44) xor data_stage(1)(46) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(56) xor data_stage(1)(62);
                crc_stage(1)(3)  <= crc_stage(0)(3) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(43) xor data_stage(1)(45) xor data_stage(1)(47) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(57) xor data_stage(1)(63);
                crc_stage(1)(4)  <= crc_stage(0)(4) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(44) xor data_stage(1)(46) xor data_stage(1)(48) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(54) xor data_stage(1)(55) xor data_stage(1)(58);
                crc_stage(1)(5)  <= crc_stage(0)(5) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(40) xor data_stage(1)(41) xor data_stage(1)(45) xor data_stage(1)(47) xor data_stage(1)(49) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(56) xor data_stage(1)(59);
                crc_stage(1)(6)  <= crc_stage(0)(6) xor data_stage(1)(33) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(41) xor data_stage(1)(44) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(56) xor data_stage(1)(57) xor data_stage(1)(62) xor data_stage(1)(63);
                crc_stage(1)(7)  <= crc_stage(0)(7) xor data_stage(1)(32) xor data_stage(1)(34) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(41) xor data_stage(1)(42) xor data_stage(1)(45) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(52) xor data_stage(1)(54) xor data_stage(1)(57) xor data_stage(1)(58) xor data_stage(1)(63);
                crc_stage(1)(8)  <= crc_stage(0)(8) xor data_stage(1)(33) xor data_stage(1)(35) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(41) xor data_stage(1)(42) xor data_stage(1)(43) xor data_stage(1)(46) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(58) xor data_stage(1)(59);
                crc_stage(1)(9)  <= crc_stage(0)(9) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(41) xor data_stage(1)(43) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(51) xor data_stage(1)(56) xor data_stage(1)(59) xor data_stage(1)(62) xor data_stage(1)(63);
                crc_stage(1)(10) <= crc_stage(0)(10) xor data_stage(1)(32) xor data_stage(1)(34) xor data_stage(1)(40) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(54) xor data_stage(1)(57) xor data_stage(1)(62);
                crc_stage(1)(11) <= crc_stage(0)(11) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(35) xor data_stage(1)(41) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(58) xor data_stage(1)(63);
                crc_stage(1)(12) <= crc_stage(0)(12) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(36) xor data_stage(1)(42) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(56) xor data_stage(1)(59);
                crc_stage(1)(13) <= crc_stage(0)(13) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(37) xor data_stage(1)(43) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(54) xor data_stage(1)(55) xor data_stage(1)(57) xor data_stage(1)(60);
                crc_stage(1)(14) <= crc_stage(0)(14) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(38) xor data_stage(1)(44) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(56) xor data_stage(1)(58) xor data_stage(1)(61);
                crc_stage(1)(15) <= crc_stage(0)(15) xor data_stage(1)(32) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(39) xor data_stage(1)(45) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(56) xor data_stage(1)(57) xor data_stage(1)(59) xor data_stage(1)(62);
                crc_stage(1)(16) <= crc_stage(0)(16) xor data_stage(1)(32) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(42) xor data_stage(1)(44) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(57) xor data_stage(1)(58) xor data_stage(1)(62);
                crc_stage(1)(17) <= crc_stage(0)(17) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(43) xor data_stage(1)(45) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(54) xor data_stage(1)(56) xor data_stage(1)(58) xor data_stage(1)(59) xor data_stage(1)(63);
                crc_stage(1)(18) <= crc_stage(0)(18) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(44) xor data_stage(1)(46) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(57) xor data_stage(1)(59) xor data_stage(1)(60);
                crc_stage(1)(19) <= crc_stage(0)(19) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(41) xor data_stage(1)(45) xor data_stage(1)(47) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(56) xor data_stage(1)(58) xor data_stage(1)(60) xor data_stage(1)(61);
                crc_stage(1)(20) <= crc_stage(0)(20) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(39) xor data_stage(1)(41) xor data_stage(1)(44) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(52) xor data_stage(1)(55) xor data_stage(1)(57) xor data_stage(1)(59) xor data_stage(1)(60) xor data_stage(1)(61) xor data_stage(1)(63);
                crc_stage(1)(21) <= crc_stage(0)(21) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(36) xor data_stage(1)(44) xor data_stage(1)(45) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(56) xor data_stage(1)(58) xor data_stage(1)(61) xor data_stage(1)(63);
                crc_stage(1)(22) <= crc_stage(0)(22) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(37) xor data_stage(1)(40) xor data_stage(1)(42) xor data_stage(1)(44) xor data_stage(1)(45) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(50) xor data_stage(1)(52) xor data_stage(1)(55) xor data_stage(1)(57) xor data_stage(1)(59) xor data_stage(1)(60) xor data_stage(1)(63);
                crc_stage(1)(23) <= crc_stage(0)(23) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(38) xor data_stage(1)(41) xor data_stage(1)(43) xor data_stage(1)(45) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(49) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(56) xor data_stage(1)(58) xor data_stage(1)(60) xor data_stage(1)(61);
                crc_stage(1)(24) <= crc_stage(0)(24) xor data_stage(1)(34) xor data_stage(1)(36) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(46) xor data_stage(1)(49) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(57) xor data_stage(1)(59) xor data_stage(1)(60) xor data_stage(1)(61) xor data_stage(1)(63);
                crc_stage(1)(25) <= crc_stage(0)(25) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(41) xor data_stage(1)(42) xor data_stage(1)(44) xor data_stage(1)(48) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(58) xor data_stage(1)(61) xor data_stage(1)(63);
                crc_stage(1)(26) <= crc_stage(0)(26) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(42) xor data_stage(1)(43) xor data_stage(1)(45) xor data_stage(1)(49) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(54) xor data_stage(1)(55) xor data_stage(1)(59) xor data_stage(1)(62);
                crc_stage(1)(27) <= crc_stage(0)(27) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(34) xor data_stage(1)(36) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(42) xor data_stage(1)(43) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(51) xor data_stage(1)(53) xor data_stage(1)(55) xor data_stage(1)(56) xor data_stage(1)(62);
                crc_stage(1)(28) <= crc_stage(0)(28) xor data_stage(1)(34) xor data_stage(1)(36) xor data_stage(1)(37) xor data_stage(1)(39) xor data_stage(1)(41) xor data_stage(1)(42) xor data_stage(1)(43) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(56) xor data_stage(1)(57) xor data_stage(1)(60) xor data_stage(1)(62);
                crc_stage(1)(29) <= crc_stage(0)(29) xor data_stage(1)(35) xor data_stage(1)(37) xor data_stage(1)(38) xor data_stage(1)(40) xor data_stage(1)(42) xor data_stage(1)(43) xor data_stage(1)(44) xor data_stage(1)(50) xor data_stage(1)(51) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(57) xor data_stage(1)(58) xor data_stage(1)(61) xor data_stage(1)(63);
                crc_stage(1)(30) <= crc_stage(0)(30) xor data_stage(1)(32) xor data_stage(1)(33) xor data_stage(1)(35) xor data_stage(1)(38) xor data_stage(1)(39) xor data_stage(1)(40) xor data_stage(1)(41) xor data_stage(1)(42) xor data_stage(1)(43) xor data_stage(1)(45) xor data_stage(1)(47) xor data_stage(1)(48) xor data_stage(1)(50) xor data_stage(1)(52) xor data_stage(1)(53) xor data_stage(1)(58) xor data_stage(1)(59) xor data_stage(1)(60) xor data_stage(1)(63);
                crc_stage(1)(31) <= crc_stage(0)(31) xor data_stage(1)(32) xor data_stage(1)(34) xor data_stage(1)(35) xor data_stage(1)(39) xor data_stage(1)(41) xor data_stage(1)(43) xor data_stage(1)(46) xor data_stage(1)(47) xor data_stage(1)(49) xor data_stage(1)(50) xor data_stage(1)(53) xor data_stage(1)(59) xor data_stage(1)(61) xor data_stage(1)(62) xor data_stage(1)(63);
            else
                crc_stage(1) <= crc_stage(0);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(2)(11 downto 8) = X"F" then
                crc_stage(2)(0)  <= crc_stage(1)(0) xor data_stage(2)(64) xor data_stage(2)(68) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(88) xor data_stage(2)(90) xor data_stage(2)(93) xor data_stage(2)(94);
                crc_stage(2)(1)  <= crc_stage(1)(1) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(69) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(79) xor data_stage(2)(80) xor data_stage(2)(89) xor data_stage(2)(91) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(2)  <= crc_stage(1)(2) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(70) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(80) xor data_stage(2)(81) xor data_stage(2)(90) xor data_stage(2)(92) xor data_stage(2)(95);
                crc_stage(2)(3)  <= crc_stage(1)(3) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(71) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(81) xor data_stage(2)(82) xor data_stage(2)(91) xor data_stage(2)(93);
                crc_stage(2)(4)  <= crc_stage(1)(4) xor data_stage(2)(64) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(68) xor data_stage(2)(72) xor data_stage(2)(79) xor data_stage(2)(80) xor data_stage(2)(82) xor data_stage(2)(83) xor data_stage(2)(92) xor data_stage(2)(94);
                crc_stage(2)(5)  <= crc_stage(1)(5) xor data_stage(2)(65) xor data_stage(2)(67) xor data_stage(2)(68) xor data_stage(2)(69) xor data_stage(2)(73) xor data_stage(2)(80) xor data_stage(2)(81) xor data_stage(2)(83) xor data_stage(2)(84) xor data_stage(2)(93) xor data_stage(2)(95);
                crc_stage(2)(6)  <= crc_stage(1)(6) xor data_stage(2)(64) xor data_stage(2)(66) xor data_stage(2)(69) xor data_stage(2)(70) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(81) xor data_stage(2)(82) xor data_stage(2)(84) xor data_stage(2)(85) xor data_stage(2)(88) xor data_stage(2)(90) xor data_stage(2)(93);
                crc_stage(2)(7)  <= crc_stage(1)(7) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(67) xor data_stage(2)(70) xor data_stage(2)(71) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(79) xor data_stage(2)(80) xor data_stage(2)(82) xor data_stage(2)(83) xor data_stage(2)(85) xor data_stage(2)(86) xor data_stage(2)(89) xor data_stage(2)(91) xor data_stage(2)(94);
                crc_stage(2)(8)  <= crc_stage(1)(8) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(68) xor data_stage(2)(71) xor data_stage(2)(72) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(80) xor data_stage(2)(81) xor data_stage(2)(83) xor data_stage(2)(84) xor data_stage(2)(86) xor data_stage(2)(87) xor data_stage(2)(90) xor data_stage(2)(92) xor data_stage(2)(95);
                crc_stage(2)(9)  <= crc_stage(1)(9) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(68) xor data_stage(2)(69) xor data_stage(2)(72) xor data_stage(2)(73) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(81) xor data_stage(2)(82) xor data_stage(2)(84) xor data_stage(2)(85) xor data_stage(2)(87) xor data_stage(2)(90) xor data_stage(2)(91) xor data_stage(2)(94);
                crc_stage(2)(10) <= crc_stage(1)(10) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(69) xor data_stage(2)(70) xor data_stage(2)(73) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(77) xor data_stage(2)(79) xor data_stage(2)(82) xor data_stage(2)(83) xor data_stage(2)(85) xor data_stage(2)(86) xor data_stage(2)(90) xor data_stage(2)(91) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(11) <= crc_stage(1)(11) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(68) xor data_stage(2)(70) xor data_stage(2)(71) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(78) xor data_stage(2)(80) xor data_stage(2)(83) xor data_stage(2)(84) xor data_stage(2)(86) xor data_stage(2)(87) xor data_stage(2)(91) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(12) <= crc_stage(1)(12) xor data_stage(2)(64) xor data_stage(2)(67) xor data_stage(2)(68) xor data_stage(2)(69) xor data_stage(2)(71) xor data_stage(2)(72) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(79) xor data_stage(2)(81) xor data_stage(2)(84) xor data_stage(2)(85) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(13) <= crc_stage(1)(13) xor data_stage(2)(65) xor data_stage(2)(68) xor data_stage(2)(69) xor data_stage(2)(70) xor data_stage(2)(72) xor data_stage(2)(73) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(80) xor data_stage(2)(82) xor data_stage(2)(85) xor data_stage(2)(86) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(14) <= crc_stage(1)(14) xor data_stage(2)(66) xor data_stage(2)(69) xor data_stage(2)(70) xor data_stage(2)(71) xor data_stage(2)(73) xor data_stage(2)(74) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(81) xor data_stage(2)(83) xor data_stage(2)(86) xor data_stage(2)(87) xor data_stage(2)(89) xor data_stage(2)(90) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(15) <= crc_stage(1)(15) xor data_stage(2)(67) xor data_stage(2)(70) xor data_stage(2)(71) xor data_stage(2)(72) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(80) xor data_stage(2)(82) xor data_stage(2)(84) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(90) xor data_stage(2)(91) xor data_stage(2)(95);
                crc_stage(2)(16) <= crc_stage(1)(16) xor data_stage(2)(64) xor data_stage(2)(71) xor data_stage(2)(72) xor data_stage(2)(73) xor data_stage(2)(78) xor data_stage(2)(80) xor data_stage(2)(81) xor data_stage(2)(83) xor data_stage(2)(85) xor data_stage(2)(89) xor data_stage(2)(90) xor data_stage(2)(91) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94);
                crc_stage(2)(17) <= crc_stage(1)(17) xor data_stage(2)(65) xor data_stage(2)(72) xor data_stage(2)(73) xor data_stage(2)(74) xor data_stage(2)(79) xor data_stage(2)(81) xor data_stage(2)(82) xor data_stage(2)(84) xor data_stage(2)(86) xor data_stage(2)(90) xor data_stage(2)(91) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(18) <= crc_stage(1)(18) xor data_stage(2)(64) xor data_stage(2)(66) xor data_stage(2)(73) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(80) xor data_stage(2)(82) xor data_stage(2)(83) xor data_stage(2)(85) xor data_stage(2)(87) xor data_stage(2)(91) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(19) <= crc_stage(1)(19) xor data_stage(2)(65) xor data_stage(2)(67) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(81) xor data_stage(2)(83) xor data_stage(2)(84) xor data_stage(2)(86) xor data_stage(2)(88) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(20) <= crc_stage(1)(20) xor data_stage(2)(64) xor data_stage(2)(66) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(82) xor data_stage(2)(84) xor data_stage(2)(85) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(90) xor data_stage(2)(95);
                crc_stage(2)(21) <= crc_stage(1)(21) xor data_stage(2)(65) xor data_stage(2)(67) xor data_stage(2)(68) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(80) xor data_stage(2)(83) xor data_stage(2)(85) xor data_stage(2)(86) xor data_stage(2)(89) xor data_stage(2)(91) xor data_stage(2)(93) xor data_stage(2)(94);
                crc_stage(2)(22) <= crc_stage(1)(22) xor data_stage(2)(66) xor data_stage(2)(69) xor data_stage(2)(75) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(81) xor data_stage(2)(84) xor data_stage(2)(86) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(95);
                crc_stage(2)(23) <= crc_stage(1)(23) xor data_stage(2)(64) xor data_stage(2)(67) xor data_stage(2)(70) xor data_stage(2)(76) xor data_stage(2)(78) xor data_stage(2)(79) xor data_stage(2)(80) xor data_stage(2)(82) xor data_stage(2)(85) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(93) xor data_stage(2)(94);
                crc_stage(2)(24) <= crc_stage(1)(24) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(71) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(80) xor data_stage(2)(81) xor data_stage(2)(83) xor data_stage(2)(86) xor data_stage(2)(89) xor data_stage(2)(93) xor data_stage(2)(95);
                crc_stage(2)(25) <= crc_stage(1)(25) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(68) xor data_stage(2)(72) xor data_stage(2)(75) xor data_stage(2)(77) xor data_stage(2)(81) xor data_stage(2)(82) xor data_stage(2)(84) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(93);
                crc_stage(2)(26) <= crc_stage(1)(26) xor data_stage(2)(64) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(69) xor data_stage(2)(73) xor data_stage(2)(76) xor data_stage(2)(78) xor data_stage(2)(82) xor data_stage(2)(83) xor data_stage(2)(85) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(94);
                crc_stage(2)(27) <= crc_stage(1)(27) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(67) xor data_stage(2)(70) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(83) xor data_stage(2)(84) xor data_stage(2)(86) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(28) <= crc_stage(1)(28) xor data_stage(2)(64) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(71) xor data_stage(2)(77) xor data_stage(2)(84) xor data_stage(2)(85) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(93) xor data_stage(2)(95);
                crc_stage(2)(29) <= crc_stage(1)(29) xor data_stage(2)(65) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(72) xor data_stage(2)(78) xor data_stage(2)(85) xor data_stage(2)(86) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(90) xor data_stage(2)(94);
                crc_stage(2)(30) <= crc_stage(1)(30) xor data_stage(2)(66) xor data_stage(2)(67) xor data_stage(2)(73) xor data_stage(2)(75) xor data_stage(2)(76) xor data_stage(2)(78) xor data_stage(2)(86) xor data_stage(2)(87) xor data_stage(2)(88) xor data_stage(2)(89) xor data_stage(2)(91) xor data_stage(2)(93) xor data_stage(2)(94) xor data_stage(2)(95);
                crc_stage(2)(31) <= crc_stage(1)(31) xor data_stage(2)(67) xor data_stage(2)(74) xor data_stage(2)(75) xor data_stage(2)(77) xor data_stage(2)(78) xor data_stage(2)(87) xor data_stage(2)(89) xor data_stage(2)(92) xor data_stage(2)(93) xor data_stage(2)(95);
            else
                crc_stage(2) <= crc_stage(1);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(3)(15 downto 12) = X"F" then
                crc_stage(3)(0)  <= crc_stage(2)(0) xor data_stage(3)(96) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(116) xor data_stage(3)(119) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126);
                crc_stage(3)(1)  <= crc_stage(2)(1) xor data_stage(3)(97) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(117) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(2)  <= crc_stage(2)(2) xor data_stage(3)(96) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(118) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(3)  <= crc_stage(2)(3) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(103) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(117) xor data_stage(3)(119) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(127);
                crc_stage(3)(4)  <= crc_stage(2)(4) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(104) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(116) xor data_stage(3)(117) xor data_stage(3)(118) xor data_stage(3)(120) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126);
                crc_stage(3)(5)  <= crc_stage(2)(5) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(103) xor data_stage(3)(105) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(117) xor data_stage(3)(118) xor data_stage(3)(119) xor data_stage(3)(121) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(6)  <= crc_stage(2)(6) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(116) xor data_stage(3)(118) xor data_stage(3)(121) xor data_stage(3)(124) xor data_stage(3)(127);
                crc_stage(3)(7)  <= crc_stage(2)(7) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(117) xor data_stage(3)(119) xor data_stage(3)(122) xor data_stage(3)(125);
                crc_stage(3)(8)  <= crc_stage(2)(8) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(118) xor data_stage(3)(120) xor data_stage(3)(123) xor data_stage(3)(126);
                crc_stage(3)(9)  <= crc_stage(2)(9) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(120) xor data_stage(3)(122) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(10) <= crc_stage(2)(10) xor data_stage(3)(96) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(117) xor data_stage(3)(119) xor data_stage(3)(120) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(127);
                crc_stage(3)(11) <= crc_stage(2)(11) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(118) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126);
                crc_stage(3)(12) <= crc_stage(2)(12) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(119) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(13) <= crc_stage(2)(13) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(116) xor data_stage(3)(117) xor data_stage(3)(120) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(14) <= crc_stage(2)(14) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(117) xor data_stage(3)(118) xor data_stage(3)(121) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(15) <= crc_stage(2)(15) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(118) xor data_stage(3)(119) xor data_stage(3)(122) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(127);
                crc_stage(3)(16) <= crc_stage(2)(16) xor data_stage(3)(97) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(106) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(117) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124);
                crc_stage(3)(17) <= crc_stage(2)(17) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(107) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(118) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125);
                crc_stage(3)(18) <= crc_stage(2)(18) xor data_stage(3)(96) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(108) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(119) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126);
                crc_stage(3)(19) <= crc_stage(2)(19) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(109) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(117) xor data_stage(3)(120) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(20) <= crc_stage(2)(20) xor data_stage(3)(97) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(104) xor data_stage(3)(106) xor data_stage(3)(108) xor data_stage(3)(110) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(117) xor data_stage(3)(118) xor data_stage(3)(119) xor data_stage(3)(120) xor data_stage(3)(122) xor data_stage(3)(124) xor data_stage(3)(127);
                crc_stage(3)(21) <= crc_stage(2)(21) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(118) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(126);
                crc_stage(3)(22) <= crc_stage(2)(22) xor data_stage(3)(96) xor data_stage(3)(98) xor data_stage(3)(100) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(114) xor data_stage(3)(117) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(23) <= crc_stage(2)(23) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(115) xor data_stage(3)(118) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(127);
                crc_stage(3)(24) <= crc_stage(2)(24) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(102) xor data_stage(3)(105) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(123) xor data_stage(3)(126);
                crc_stage(3)(25) <= crc_stage(2)(25) xor data_stage(3)(97) xor data_stage(3)(100) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(109) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(113) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(119) xor data_stage(3)(120) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(26) <= crc_stage(2)(26) xor data_stage(3)(98) xor data_stage(3)(101) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(108) xor data_stage(3)(110) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(114) xor data_stage(3)(116) xor data_stage(3)(117) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(27) <= crc_stage(2)(27) xor data_stage(3)(96) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(106) xor data_stage(3)(109) xor data_stage(3)(111) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(117) xor data_stage(3)(118) xor data_stage(3)(119) xor data_stage(3)(120) xor data_stage(3)(124) xor data_stage(3)(125) xor data_stage(3)(126) xor data_stage(3)(127);
                crc_stage(3)(28) <= crc_stage(2)(28) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(106) xor data_stage(3)(108) xor data_stage(3)(110) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(117) xor data_stage(3)(118) xor data_stage(3)(122) xor data_stage(3)(124) xor data_stage(3)(127);
                crc_stage(3)(29) <= crc_stage(2)(29) xor data_stage(3)(96) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(100) xor data_stage(3)(102) xor data_stage(3)(107) xor data_stage(3)(109) xor data_stage(3)(111) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(116) xor data_stage(3)(118) xor data_stage(3)(119) xor data_stage(3)(123) xor data_stage(3)(125);
                crc_stage(3)(30) <= crc_stage(2)(30) xor data_stage(3)(96) xor data_stage(3)(97) xor data_stage(3)(98) xor data_stage(3)(99) xor data_stage(3)(101) xor data_stage(3)(104) xor data_stage(3)(105) xor data_stage(3)(107) xor data_stage(3)(110) xor data_stage(3)(113) xor data_stage(3)(114) xor data_stage(3)(115) xor data_stage(3)(117) xor data_stage(3)(121) xor data_stage(3)(122) xor data_stage(3)(125);
                crc_stage(3)(31) <= crc_stage(2)(31) xor data_stage(3)(97) xor data_stage(3)(99) xor data_stage(3)(102) xor data_stage(3)(103) xor data_stage(3)(104) xor data_stage(3)(106) xor data_stage(3)(107) xor data_stage(3)(111) xor data_stage(3)(112) xor data_stage(3)(113) xor data_stage(3)(115) xor data_stage(3)(118) xor data_stage(3)(119) xor data_stage(3)(120) xor data_stage(3)(121) xor data_stage(3)(123) xor data_stage(3)(124) xor data_stage(3)(125);
            else
                crc_stage(3) <= crc_stage(2);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(4)(19 downto 16) = X"F" then
                crc_stage(4)(0)  <= crc_stage(3)(0) xor data_stage(4)(131) xor data_stage(4)(134) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(146) xor data_stage(4)(149) xor data_stage(4)(150) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(159);
                crc_stage(4)(1)  <= crc_stage(3)(1) xor data_stage(4)(132) xor data_stage(4)(135) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(147) xor data_stage(4)(150) xor data_stage(4)(151) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(156);
                crc_stage(4)(2)  <= crc_stage(3)(2) xor data_stage(4)(128) xor data_stage(4)(133) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(142) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(148) xor data_stage(4)(151) xor data_stage(4)(152) xor data_stage(4)(155) xor data_stage(4)(156) xor data_stage(4)(157);
                crc_stage(4)(3)  <= crc_stage(3)(3) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(134) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(146) xor data_stage(4)(147) xor data_stage(4)(149) xor data_stage(4)(152) xor data_stage(4)(153) xor data_stage(4)(156) xor data_stage(4)(157) xor data_stage(4)(158);
                crc_stage(4)(4)  <= crc_stage(3)(4) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(135) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(142) xor data_stage(4)(144) xor data_stage(4)(147) xor data_stage(4)(148) xor data_stage(4)(150) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(157) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(5)  <= crc_stage(3)(5) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(136) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(145) xor data_stage(4)(148) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(6)  <= crc_stage(3)(6) xor data_stage(4)(128) xor data_stage(4)(130) xor data_stage(4)(132) xor data_stage(4)(134) xor data_stage(4)(136) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(142) xor data_stage(4)(143) xor data_stage(4)(152) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(156);
                crc_stage(4)(7)  <= crc_stage(3)(7) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(131) xor data_stage(4)(133) xor data_stage(4)(135) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(157);
                crc_stage(4)(8)  <= crc_stage(3)(8) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(132) xor data_stage(4)(134) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(140) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(156) xor data_stage(4)(158);
                crc_stage(4)(9)  <= crc_stage(3)(9) xor data_stage(4)(130) xor data_stage(4)(133) xor data_stage(4)(134) xor data_stage(4)(135) xor data_stage(4)(136) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(149) xor data_stage(4)(150) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(156) xor data_stage(4)(157);
                crc_stage(4)(10) <= crc_stage(3)(10) xor data_stage(4)(128) xor data_stage(4)(135) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(142) xor data_stage(4)(143) xor data_stage(4)(145) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(153) xor data_stage(4)(157) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(11) <= crc_stage(3)(11) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(146) xor data_stage(4)(150) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(12) <= crc_stage(3)(12) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(147) xor data_stage(4)(151) xor data_stage(4)(153) xor data_stage(4)(155) xor data_stage(4)(159);
                crc_stage(4)(13) <= crc_stage(3)(13) xor data_stage(4)(128) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(142) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(148) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(156);
                crc_stage(4)(14) <= crc_stage(3)(14) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(146) xor data_stage(4)(147) xor data_stage(4)(149) xor data_stage(4)(153) xor data_stage(4)(155) xor data_stage(4)(157);
                crc_stage(4)(15) <= crc_stage(3)(15) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(140) xor data_stage(4)(142) xor data_stage(4)(144) xor data_stage(4)(147) xor data_stage(4)(148) xor data_stage(4)(150) xor data_stage(4)(154) xor data_stage(4)(156) xor data_stage(4)(158);
                crc_stage(4)(16) <= crc_stage(3)(16) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(133) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(141) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(148) xor data_stage(4)(150) xor data_stage(4)(151) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(157);
                crc_stage(4)(17) <= crc_stage(3)(17) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(134) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(142) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(147) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(158);
                crc_stage(4)(18) <= crc_stage(3)(18) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(135) xor data_stage(4)(138) xor data_stage(4)(140) xor data_stage(4)(142) xor data_stage(4)(143) xor data_stage(4)(146) xor data_stage(4)(147) xor data_stage(4)(148) xor data_stage(4)(150) xor data_stage(4)(152) xor data_stage(4)(153) xor data_stage(4)(155) xor data_stage(4)(156) xor data_stage(4)(159);
                crc_stage(4)(19) <= crc_stage(3)(19) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(136) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(147) xor data_stage(4)(148) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(156) xor data_stage(4)(157);
                crc_stage(4)(20) <= crc_stage(3)(20) xor data_stage(4)(128) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(136) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(142) xor data_stage(4)(143) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(148) xor data_stage(4)(152) xor data_stage(4)(153) xor data_stage(4)(157) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(21) <= crc_stage(3)(21) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(136) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(140) xor data_stage(4)(147) xor data_stage(4)(150) xor data_stage(4)(155) xor data_stage(4)(158);
                crc_stage(4)(22) <= crc_stage(3)(22) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(136) xor data_stage(4)(137) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(146) xor data_stage(4)(148) xor data_stage(4)(149) xor data_stage(4)(150) xor data_stage(4)(151) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(156);
                crc_stage(4)(23) <= crc_stage(3)(23) xor data_stage(4)(128) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(134) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(142) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(147) xor data_stage(4)(149) xor data_stage(4)(150) xor data_stage(4)(151) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(155) xor data_stage(4)(156) xor data_stage(4)(157);
                crc_stage(4)(24) <= crc_stage(3)(24) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(135) xor data_stage(4)(136) xor data_stage(4)(139) xor data_stage(4)(140) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(148) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(156) xor data_stage(4)(157) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(25) <= crc_stage(3)(25) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(133) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(157) xor data_stage(4)(158);
                crc_stage(4)(26) <= crc_stage(3)(26) xor data_stage(4)(128) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(134) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(142) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(153) xor data_stage(4)(155) xor data_stage(4)(158) xor data_stage(4)(159);
                crc_stage(4)(27) <= crc_stage(3)(27) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(134) xor data_stage(4)(135) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(147) xor data_stage(4)(149) xor data_stage(4)(150) xor data_stage(4)(153) xor data_stage(4)(155) xor data_stage(4)(156);
                crc_stage(4)(28) <= crc_stage(3)(28) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(133) xor data_stage(4)(135) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(148) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(153) xor data_stage(4)(155) xor data_stage(4)(156) xor data_stage(4)(157) xor data_stage(4)(159);
                crc_stage(4)(29) <= crc_stage(3)(29) xor data_stage(4)(128) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(131) xor data_stage(4)(132) xor data_stage(4)(134) xor data_stage(4)(136) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(140) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(146) xor data_stage(4)(149) xor data_stage(4)(150) xor data_stage(4)(152) xor data_stage(4)(154) xor data_stage(4)(156) xor data_stage(4)(157) xor data_stage(4)(158);
                crc_stage(4)(30) <= crc_stage(3)(30) xor data_stage(4)(129) xor data_stage(4)(130) xor data_stage(4)(132) xor data_stage(4)(133) xor data_stage(4)(134) xor data_stage(4)(135) xor data_stage(4)(136) xor data_stage(4)(137) xor data_stage(4)(138) xor data_stage(4)(139) xor data_stage(4)(141) xor data_stage(4)(143) xor data_stage(4)(144) xor data_stage(4)(145) xor data_stage(4)(147) xor data_stage(4)(149) xor data_stage(4)(151) xor data_stage(4)(154) xor data_stage(4)(157) xor data_stage(4)(158);
                crc_stage(4)(31) <= crc_stage(3)(31) xor data_stage(4)(130) xor data_stage(4)(133) xor data_stage(4)(135) xor data_stage(4)(137) xor data_stage(4)(139) xor data_stage(4)(142) xor data_stage(4)(143) xor data_stage(4)(145) xor data_stage(4)(148) xor data_stage(4)(149) xor data_stage(4)(152) xor data_stage(4)(153) xor data_stage(4)(154) xor data_stage(4)(158);
            else
                crc_stage(4) <= crc_stage(3);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(5)(23 downto 20) = X"F" then
                crc_stage(5)(0)  <= crc_stage(4)(0) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(184) xor data_stage(5)(185) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(1)  <= crc_stage(4)(1) xor data_stage(5)(160) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(171) xor data_stage(5)(172) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(191);
                crc_stage(5)(2)  <= crc_stage(4)(2) xor data_stage(5)(161) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(177) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(186) xor data_stage(5)(187);
                crc_stage(5)(3)  <= crc_stage(4)(3) xor data_stage(5)(162) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(176) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(187) xor data_stage(5)(188);
                crc_stage(5)(4)  <= crc_stage(4)(4) xor data_stage(5)(163) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(171) xor data_stage(5)(172) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(188) xor data_stage(5)(189);
                crc_stage(5)(5)  <= crc_stage(4)(5) xor data_stage(5)(160) xor data_stage(5)(164) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(184) xor data_stage(5)(189) xor data_stage(5)(190);
                crc_stage(5)(6)  <= crc_stage(4)(6) xor data_stage(5)(160) xor data_stage(5)(161) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(183);
                crc_stage(5)(7)  <= crc_stage(4)(7) xor data_stage(5)(161) xor data_stage(5)(162) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(176) xor data_stage(5)(177) xor data_stage(5)(179) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(184);
                crc_stage(5)(8)  <= crc_stage(4)(8) xor data_stage(5)(162) xor data_stage(5)(163) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(180) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(185);
                crc_stage(5)(9)  <= crc_stage(4)(9) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(168) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(177) xor data_stage(5)(181) xor data_stage(5)(183) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(10) <= crc_stage(4)(10) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(176) xor data_stage(5)(177) xor data_stage(5)(179) xor data_stage(5)(182) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(187) xor data_stage(5)(190);
                crc_stage(5)(11) <= crc_stage(4)(11) xor data_stage(5)(160) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(172) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(180) xor data_stage(5)(183) xor data_stage(5)(186) xor data_stage(5)(187) xor data_stage(5)(188) xor data_stage(5)(191);
                crc_stage(5)(12) <= crc_stage(4)(12) xor data_stage(5)(160) xor data_stage(5)(161) xor data_stage(5)(165) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(181) xor data_stage(5)(184) xor data_stage(5)(187) xor data_stage(5)(188) xor data_stage(5)(189);
                crc_stage(5)(13) <= crc_stage(4)(13) xor data_stage(5)(160) xor data_stage(5)(161) xor data_stage(5)(162) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(171) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(182) xor data_stage(5)(185) xor data_stage(5)(188) xor data_stage(5)(189) xor data_stage(5)(190);
                crc_stage(5)(14) <= crc_stage(4)(14) xor data_stage(5)(161) xor data_stage(5)(162) xor data_stage(5)(163) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(183) xor data_stage(5)(186) xor data_stage(5)(189) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(15) <= crc_stage(4)(15) xor data_stage(5)(162) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(184) xor data_stage(5)(187) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(16) <= crc_stage(4)(16) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(184) xor data_stage(5)(188) xor data_stage(5)(190);
                crc_stage(5)(17) <= crc_stage(4)(17) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(177) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(183) xor data_stage(5)(184) xor data_stage(5)(185) xor data_stage(5)(189) xor data_stage(5)(191);
                crc_stage(5)(18) <= crc_stage(4)(18) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(178) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(184) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(190);
                crc_stage(5)(19) <= crc_stage(4)(19) xor data_stage(5)(160) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(172) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(179) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(187) xor data_stage(5)(191);
                crc_stage(5)(20) <= crc_stage(4)(20) xor data_stage(5)(161) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(170) xor data_stage(5)(172) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(184) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(187) xor data_stage(5)(188) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(21) <= crc_stage(4)(21) xor data_stage(5)(160) xor data_stage(5)(162) xor data_stage(5)(163) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(174) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(183) xor data_stage(5)(186) xor data_stage(5)(187) xor data_stage(5)(188) xor data_stage(5)(189) xor data_stage(5)(190);
                crc_stage(5)(22) <= crc_stage(4)(22) xor data_stage(5)(161) xor data_stage(5)(165) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(178) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(185) xor data_stage(5)(187) xor data_stage(5)(188) xor data_stage(5)(189);
                crc_stage(5)(23) <= crc_stage(4)(23) xor data_stage(5)(162) xor data_stage(5)(166) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(179) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(186) xor data_stage(5)(188) xor data_stage(5)(189) xor data_stage(5)(190);
                crc_stage(5)(24) <= crc_stage(4)(24) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(168) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(176) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(180) xor data_stage(5)(183) xor data_stage(5)(185) xor data_stage(5)(187) xor data_stage(5)(189);
                crc_stage(5)(25) <= crc_stage(4)(25) xor data_stage(5)(160) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(180) xor data_stage(5)(181) xor data_stage(5)(185) xor data_stage(5)(186) xor data_stage(5)(188) xor data_stage(5)(191);
                crc_stage(5)(26) <= crc_stage(4)(26) xor data_stage(5)(161) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(181) xor data_stage(5)(182) xor data_stage(5)(186) xor data_stage(5)(187) xor data_stage(5)(189);
                crc_stage(5)(27) <= crc_stage(4)(27) xor data_stage(5)(160) xor data_stage(5)(162) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(169) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(179) xor data_stage(5)(182) xor data_stage(5)(183) xor data_stage(5)(184) xor data_stage(5)(185) xor data_stage(5)(187) xor data_stage(5)(188) xor data_stage(5)(191);
                crc_stage(5)(28) <= crc_stage(4)(28) xor data_stage(5)(161) xor data_stage(5)(171) xor data_stage(5)(175) xor data_stage(5)(177) xor data_stage(5)(180) xor data_stage(5)(183) xor data_stage(5)(186) xor data_stage(5)(188) xor data_stage(5)(189) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(29) <= crc_stage(4)(29) xor data_stage(5)(160) xor data_stage(5)(162) xor data_stage(5)(172) xor data_stage(5)(176) xor data_stage(5)(178) xor data_stage(5)(181) xor data_stage(5)(184) xor data_stage(5)(187) xor data_stage(5)(189) xor data_stage(5)(190) xor data_stage(5)(191);
                crc_stage(5)(30) <= crc_stage(4)(30) xor data_stage(5)(161) xor data_stage(5)(164) xor data_stage(5)(165) xor data_stage(5)(167) xor data_stage(5)(168) xor data_stage(5)(170) xor data_stage(5)(171) xor data_stage(5)(174) xor data_stage(5)(175) xor data_stage(5)(178) xor data_stage(5)(182) xor data_stage(5)(184) xor data_stage(5)(188);
                crc_stage(5)(31) <= crc_stage(4)(31) xor data_stage(5)(162) xor data_stage(5)(163) xor data_stage(5)(164) xor data_stage(5)(166) xor data_stage(5)(167) xor data_stage(5)(169) xor data_stage(5)(170) xor data_stage(5)(172) xor data_stage(5)(173) xor data_stage(5)(174) xor data_stage(5)(176) xor data_stage(5)(177) xor data_stage(5)(178) xor data_stage(5)(183) xor data_stage(5)(184) xor data_stage(5)(189) xor data_stage(5)(190) xor data_stage(5)(191);
            else
                crc_stage(5) <= crc_stage(4);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(6)(27 downto 24) = X"F" then
                crc_stage(6)(0)  <= crc_stage(5)(0) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(197) xor data_stage(6)(200) xor data_stage(6)(202) xor data_stage(6)(203) xor data_stage(6)(207) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(222);
                crc_stage(6)(1)  <= crc_stage(5)(1) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(198) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(208) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(2)  <= crc_stage(5)(2) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(199) xor data_stage(6)(202) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(209) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(222);
                crc_stage(6)(3)  <= crc_stage(5)(3) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(200) xor data_stage(6)(203) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(210) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(4)  <= crc_stage(5)(4) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(201) xor data_stage(6)(204) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(211) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(221) xor data_stage(6)(222);
                crc_stage(6)(5)  <= crc_stage(5)(5) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(202) xor data_stage(6)(205) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(212) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(221) xor data_stage(6)(222) xor data_stage(6)(223);
                crc_stage(6)(6)  <= crc_stage(5)(6) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(201) xor data_stage(6)(202) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(210) xor data_stage(6)(212) xor data_stage(6)(214) xor data_stage(6)(217) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(7)  <= crc_stage(5)(7) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(202) xor data_stage(6)(203) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(211) xor data_stage(6)(213) xor data_stage(6)(215) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(222);
                crc_stage(6)(8)  <= crc_stage(5)(8) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(200) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(212) xor data_stage(6)(214) xor data_stage(6)(216) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(9)  <= crc_stage(5)(9) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(196) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(207) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(214) xor data_stage(6)(216) xor data_stage(6)(218);
                crc_stage(6)(10) <= crc_stage(5)(10) xor data_stage(6)(199) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(214) xor data_stage(6)(216) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(222);
                crc_stage(6)(11) <= crc_stage(5)(11) xor data_stage(6)(200) xor data_stage(6)(202) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(215) xor data_stage(6)(217) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(12) <= crc_stage(5)(12) xor data_stage(6)(192) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(216) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(221) xor data_stage(6)(222);
                crc_stage(6)(13) <= crc_stage(5)(13) xor data_stage(6)(193) xor data_stage(6)(202) xor data_stage(6)(204) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(217) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(222) xor data_stage(6)(223);
                crc_stage(6)(14) <= crc_stage(5)(14) xor data_stage(6)(194) xor data_stage(6)(203) xor data_stage(6)(205) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(222) xor data_stage(6)(223);
                crc_stage(6)(15) <= crc_stage(5)(15) xor data_stage(6)(192) xor data_stage(6)(195) xor data_stage(6)(204) xor data_stage(6)(206) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(16) <= crc_stage(5)(16) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(200) xor data_stage(6)(202) xor data_stage(6)(203) xor data_stage(6)(205) xor data_stage(6)(211) xor data_stage(6)(217) xor data_stage(6)(218);
                crc_stage(6)(17) <= crc_stage(5)(17) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(206) xor data_stage(6)(212) xor data_stage(6)(218) xor data_stage(6)(219);
                crc_stage(6)(18) <= crc_stage(5)(18) xor data_stage(6)(192) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(202) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(207) xor data_stage(6)(213) xor data_stage(6)(219) xor data_stage(6)(220);
                crc_stage(6)(19) <= crc_stage(5)(19) xor data_stage(6)(193) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(203) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(208) xor data_stage(6)(214) xor data_stage(6)(220) xor data_stage(6)(221);
                crc_stage(6)(20) <= crc_stage(5)(20) xor data_stage(6)(193) xor data_stage(6)(195) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(201) xor data_stage(6)(202) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(206) xor data_stage(6)(210) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(221);
                crc_stage(6)(21) <= crc_stage(5)(21) xor data_stage(6)(193) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(216) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(221);
                crc_stage(6)(22) <= crc_stage(5)(22) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(202) xor data_stage(6)(203) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(209) xor data_stage(6)(211) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(218) xor data_stage(6)(221);
                crc_stage(6)(23) <= crc_stage(5)(23) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(210) xor data_stage(6)(212) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(219) xor data_stage(6)(222);
                crc_stage(6)(24) <= crc_stage(5)(24) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(198) xor data_stage(6)(201) xor data_stage(6)(202) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(208) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(222) xor data_stage(6)(223);
                crc_stage(6)(25) <= crc_stage(5)(25) xor data_stage(6)(192) xor data_stage(6)(195) xor data_stage(6)(197) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(214) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(222) xor data_stage(6)(223);
                crc_stage(6)(26) <= crc_stage(5)(26) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(196) xor data_stage(6)(198) xor data_stage(6)(200) xor data_stage(6)(201) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(208) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(215) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(223);
                crc_stage(6)(27) <= crc_stage(5)(27) xor data_stage(6)(192) xor data_stage(6)(195) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(206) xor data_stage(6)(208) xor data_stage(6)(210) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219);
                crc_stage(6)(28) <= crc_stage(5)(28) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(201) xor data_stage(6)(203) xor data_stage(6)(204) xor data_stage(6)(210) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(217) xor data_stage(6)(219) xor data_stage(6)(222);
                crc_stage(6)(29) <= crc_stage(5)(29) xor data_stage(6)(192) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(197) xor data_stage(6)(198) xor data_stage(6)(202) xor data_stage(6)(204) xor data_stage(6)(205) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(218) xor data_stage(6)(220) xor data_stage(6)(223);
                crc_stage(6)(30) <= crc_stage(5)(30) xor data_stage(6)(194) xor data_stage(6)(195) xor data_stage(6)(196) xor data_stage(6)(198) xor data_stage(6)(199) xor data_stage(6)(200) xor data_stage(6)(202) xor data_stage(6)(205) xor data_stage(6)(206) xor data_stage(6)(207) xor data_stage(6)(209) xor data_stage(6)(210) xor data_stage(6)(217) xor data_stage(6)(218) xor data_stage(6)(219) xor data_stage(6)(220) xor data_stage(6)(221) xor data_stage(6)(222);
                crc_stage(6)(31) <= crc_stage(5)(31) xor data_stage(6)(192) xor data_stage(6)(193) xor data_stage(6)(194) xor data_stage(6)(196) xor data_stage(6)(199) xor data_stage(6)(201) xor data_stage(6)(202) xor data_stage(6)(206) xor data_stage(6)(208) xor data_stage(6)(209) xor data_stage(6)(211) xor data_stage(6)(212) xor data_stage(6)(213) xor data_stage(6)(214) xor data_stage(6)(215) xor data_stage(6)(216) xor data_stage(6)(217) xor data_stage(6)(219) xor data_stage(6)(221) xor data_stage(6)(223);
            else
                crc_stage(6) <= crc_stage(5);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(7)(31 downto 28) = X"F" then
                crc_stage(7)(0)  <= crc_stage(6)(0) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(226) xor data_stage(7)(229) xor data_stage(7)(233) xor data_stage(7)(235) xor data_stage(7)(236) xor data_stage(7)(238) xor data_stage(7)(239) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(251) xor data_stage(7)(253) xor data_stage(7)(255);
                crc_stage(7)(1)  <= crc_stage(6)(1) xor data_stage(7)(225) xor data_stage(7)(226) xor data_stage(7)(227) xor data_stage(7)(230) xor data_stage(7)(234) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(240) xor data_stage(7)(244) xor data_stage(7)(245) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(252) xor data_stage(7)(254);
                crc_stage(7)(2)  <= crc_stage(6)(2) xor data_stage(7)(224) xor data_stage(7)(226) xor data_stage(7)(227) xor data_stage(7)(228) xor data_stage(7)(231) xor data_stage(7)(235) xor data_stage(7)(237) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(241) xor data_stage(7)(245) xor data_stage(7)(246) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(253) xor data_stage(7)(255);
                crc_stage(7)(3)  <= crc_stage(6)(3) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(232) xor data_stage(7)(236) xor data_stage(7)(238) xor data_stage(7)(239) xor data_stage(7)(241) xor data_stage(7)(242) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(254);
                crc_stage(7)(4)  <= crc_stage(6)(4) xor data_stage(7)(224) xor data_stage(7)(226) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(233) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(240) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(255);
                crc_stage(7)(5)  <= crc_stage(6)(5) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(234) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(241) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(252) xor data_stage(7)(253);
                crc_stage(7)(6)  <= crc_stage(6)(6) xor data_stage(7)(225) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(236) xor data_stage(7)(238) xor data_stage(7)(241) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(245) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(7)  <= crc_stage(6)(7) xor data_stage(7)(224) xor data_stage(7)(226) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(234) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(246) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(255);
                crc_stage(7)(8)  <= crc_stage(6)(8) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(234) xor data_stage(7)(235) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(245) xor data_stage(7)(247) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(253);
                crc_stage(7)(9)  <= crc_stage(6)(9) xor data_stage(7)(225) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(238) xor data_stage(7)(241) xor data_stage(7)(243) xor data_stage(7)(245) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(250) xor data_stage(7)(252) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(10) <= crc_stage(6)(10) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(230) xor data_stage(7)(232) xor data_stage(7)(236) xor data_stage(7)(238) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(246);
                crc_stage(7)(11) <= crc_stage(6)(11) xor data_stage(7)(225) xor data_stage(7)(226) xor data_stage(7)(231) xor data_stage(7)(233) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(247);
                crc_stage(7)(12) <= crc_stage(6)(12) xor data_stage(7)(224) xor data_stage(7)(226) xor data_stage(7)(227) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(244) xor data_stage(7)(245) xor data_stage(7)(248);
                crc_stage(7)(13) <= crc_stage(6)(13) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(228) xor data_stage(7)(233) xor data_stage(7)(235) xor data_stage(7)(239) xor data_stage(7)(241) xor data_stage(7)(245) xor data_stage(7)(246) xor data_stage(7)(249);
                crc_stage(7)(14) <= crc_stage(6)(14) xor data_stage(7)(224) xor data_stage(7)(226) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(234) xor data_stage(7)(236) xor data_stage(7)(240) xor data_stage(7)(242) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(250);
                crc_stage(7)(15) <= crc_stage(6)(15) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(235) xor data_stage(7)(237) xor data_stage(7)(241) xor data_stage(7)(243) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(251);
                crc_stage(7)(16) <= crc_stage(6)(16) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(233) xor data_stage(7)(235) xor data_stage(7)(239) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(247) xor data_stage(7)(249) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(253) xor data_stage(7)(255);
                crc_stage(7)(17) <= crc_stage(6)(17) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(236) xor data_stage(7)(240) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(248) xor data_stage(7)(250) xor data_stage(7)(252) xor data_stage(7)(253) xor data_stage(7)(254);
                crc_stage(7)(18) <= crc_stage(6)(18) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(235) xor data_stage(7)(237) xor data_stage(7)(241) xor data_stage(7)(244) xor data_stage(7)(245) xor data_stage(7)(249) xor data_stage(7)(251) xor data_stage(7)(253) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(19) <= crc_stage(6)(19) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(234) xor data_stage(7)(236) xor data_stage(7)(238) xor data_stage(7)(242) xor data_stage(7)(245) xor data_stage(7)(246) xor data_stage(7)(250) xor data_stage(7)(252) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(20) <= crc_stage(6)(20) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(226) xor data_stage(7)(229) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(238) xor data_stage(7)(244) xor data_stage(7)(246) xor data_stage(7)(248);
                crc_stage(7)(21) <= crc_stage(6)(21) xor data_stage(7)(224) xor data_stage(7)(227) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(245) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(251) xor data_stage(7)(253) xor data_stage(7)(255);
                crc_stage(7)(22) <= crc_stage(6)(22) xor data_stage(7)(224) xor data_stage(7)(226) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(233) xor data_stage(7)(235) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(243) xor data_stage(7)(245) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(253) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(23) <= crc_stage(6)(23) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(244) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(253) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(24) <= crc_stage(6)(24) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(228) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(241) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(245) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(252) xor data_stage(7)(254);
                crc_stage(7)(25) <= crc_stage(6)(25) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(235) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(245) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(250);
                crc_stage(7)(26) <= crc_stage(6)(26) xor data_stage(7)(224) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(251);
                crc_stage(7)(27) <= crc_stage(6)(27) xor data_stage(7)(226) xor data_stage(7)(229) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(235) xor data_stage(7)(236) xor data_stage(7)(237) xor data_stage(7)(241) xor data_stage(7)(243) xor data_stage(7)(245) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(253) xor data_stage(7)(255);
                crc_stage(7)(28) <= crc_stage(6)(28) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(226) xor data_stage(7)(227) xor data_stage(7)(229) xor data_stage(7)(230) xor data_stage(7)(237) xor data_stage(7)(239) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(250) xor data_stage(7)(252) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(29) <= crc_stage(6)(29) xor data_stage(7)(225) xor data_stage(7)(226) xor data_stage(7)(227) xor data_stage(7)(228) xor data_stage(7)(230) xor data_stage(7)(231) xor data_stage(7)(238) xor data_stage(7)(240) xor data_stage(7)(243) xor data_stage(7)(244) xor data_stage(7)(247) xor data_stage(7)(248) xor data_stage(7)(249) xor data_stage(7)(251) xor data_stage(7)(253) xor data_stage(7)(255);
                crc_stage(7)(30) <= crc_stage(6)(30) xor data_stage(7)(225) xor data_stage(7)(227) xor data_stage(7)(228) xor data_stage(7)(231) xor data_stage(7)(232) xor data_stage(7)(233) xor data_stage(7)(235) xor data_stage(7)(236) xor data_stage(7)(238) xor data_stage(7)(241) xor data_stage(7)(243) xor data_stage(7)(245) xor data_stage(7)(247) xor data_stage(7)(249) xor data_stage(7)(250) xor data_stage(7)(251) xor data_stage(7)(252) xor data_stage(7)(253) xor data_stage(7)(254) xor data_stage(7)(255);
                crc_stage(7)(31) <= crc_stage(6)(31) xor data_stage(7)(224) xor data_stage(7)(225) xor data_stage(7)(228) xor data_stage(7)(232) xor data_stage(7)(234) xor data_stage(7)(235) xor data_stage(7)(237) xor data_stage(7)(238) xor data_stage(7)(242) xor data_stage(7)(243) xor data_stage(7)(246) xor data_stage(7)(247) xor data_stage(7)(250) xor data_stage(7)(252) xor data_stage(7)(254);
            else
                crc_stage(8) <= crc_stage(6);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(8)(35 downto 32) = X"F" then
                crc_stage(8)(0)  <= crc_stage(7)(0) xor data_stage(8)(257) xor data_stage(8)(260) xor data_stage(8)(264) xor data_stage(8)(269) xor data_stage(8)(275) xor data_stage(8)(278) xor data_stage(8)(282) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(286);
                crc_stage(8)(1)  <= crc_stage(7)(1) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(261) xor data_stage(8)(265) xor data_stage(8)(270) xor data_stage(8)(276) xor data_stage(8)(279) xor data_stage(8)(283) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(2)  <= crc_stage(7)(2) xor data_stage(8)(257) xor data_stage(8)(259) xor data_stage(8)(262) xor data_stage(8)(266) xor data_stage(8)(271) xor data_stage(8)(277) xor data_stage(8)(280) xor data_stage(8)(284) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(3)  <= crc_stage(7)(3) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(260) xor data_stage(8)(263) xor data_stage(8)(267) xor data_stage(8)(272) xor data_stage(8)(278) xor data_stage(8)(281) xor data_stage(8)(285) xor data_stage(8)(287);
                crc_stage(8)(4)  <= crc_stage(7)(4) xor data_stage(8)(257) xor data_stage(8)(259) xor data_stage(8)(261) xor data_stage(8)(264) xor data_stage(8)(268) xor data_stage(8)(273) xor data_stage(8)(279) xor data_stage(8)(282) xor data_stage(8)(286);
                crc_stage(8)(5)  <= crc_stage(7)(5) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(265) xor data_stage(8)(269) xor data_stage(8)(274) xor data_stage(8)(280) xor data_stage(8)(283) xor data_stage(8)(287);
                crc_stage(8)(6)  <= crc_stage(7)(6) xor data_stage(8)(259) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(266) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(278) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(285) xor data_stage(8)(286);
                crc_stage(8)(7)  <= crc_stage(7)(7) xor data_stage(8)(256) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(267) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(279) xor data_stage(8)(282) xor data_stage(8)(283) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(8)  <= crc_stage(7)(8) xor data_stage(8)(256) xor data_stage(8)(257) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(268) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(280) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(287);
                crc_stage(8)(9)  <= crc_stage(7)(9) xor data_stage(8)(258) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(275) xor data_stage(8)(278) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(286);
                crc_stage(8)(10) <= crc_stage(7)(10) xor data_stage(8)(256) xor data_stage(8)(257) xor data_stage(8)(259) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(269) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(11) <= crc_stage(7)(11) xor data_stage(8)(257) xor data_stage(8)(258) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(264) xor data_stage(8)(268) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(274) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(12) <= crc_stage(7)(12) xor data_stage(8)(258) xor data_stage(8)(259) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(265) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(278) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(13) <= crc_stage(7)(13) xor data_stage(8)(259) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(266) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(14) <= crc_stage(7)(14) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(267) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(277) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(282) xor data_stage(8)(283) xor data_stage(8)(287);
                crc_stage(8)(15) <= crc_stage(7)(15) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(268) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(283) xor data_stage(8)(284);
                crc_stage(8)(16) <= crc_stage(7)(16) xor data_stage(8)(257) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(286);
                crc_stage(8)(17) <= crc_stage(7)(17) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(274) xor data_stage(8)(275) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(287);
                crc_stage(8)(18) <= crc_stage(7)(18) xor data_stage(8)(257) xor data_stage(8)(259) xor data_stage(8)(262) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(269) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(283);
                crc_stage(8)(19) <= crc_stage(7)(19) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(260) xor data_stage(8)(263) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(283) xor data_stage(8)(284);
                crc_stage(8)(20) <= crc_stage(7)(20) xor data_stage(8)(256) xor data_stage(8)(259) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(275) xor data_stage(8)(277) xor data_stage(8)(283) xor data_stage(8)(286);
                crc_stage(8)(21) <= crc_stage(7)(21) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(264) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(282) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(22) <= crc_stage(7)(22) xor data_stage(8)(256) xor data_stage(8)(257) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(268) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(278) xor data_stage(8)(282) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(287);
                crc_stage(8)(23) <= crc_stage(7)(23) xor data_stage(8)(256) xor data_stage(8)(257) xor data_stage(8)(258) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(269) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(286);
                crc_stage(8)(24) <= crc_stage(7)(24) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(259) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(274) xor data_stage(8)(277) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(282) xor data_stage(8)(287);
                crc_stage(8)(25) <= crc_stage(7)(25) xor data_stage(8)(259) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(286);
                crc_stage(8)(26) <= crc_stage(7)(26) xor data_stage(8)(260) xor data_stage(8)(262) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(269) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(27) <= crc_stage(7)(27) xor data_stage(8)(257) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(263) xor data_stage(8)(264) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(268) xor data_stage(8)(270) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(275) xor data_stage(8)(278) xor data_stage(8)(283) xor data_stage(8)(287);
                crc_stage(8)(28) <= crc_stage(7)(28) xor data_stage(8)(256) xor data_stage(8)(257) xor data_stage(8)(258) xor data_stage(8)(260) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(265) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(271) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(278) xor data_stage(8)(279) xor data_stage(8)(282) xor data_stage(8)(285) xor data_stage(8)(286);
                crc_stage(8)(29) <= crc_stage(7)(29) xor data_stage(8)(256) xor data_stage(8)(257) xor data_stage(8)(258) xor data_stage(8)(259) xor data_stage(8)(261) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(266) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(272) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(275) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(279) xor data_stage(8)(280) xor data_stage(8)(283) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(30) <= crc_stage(7)(30) xor data_stage(8)(256) xor data_stage(8)(258) xor data_stage(8)(259) xor data_stage(8)(262) xor data_stage(8)(263) xor data_stage(8)(267) xor data_stage(8)(268) xor data_stage(8)(273) xor data_stage(8)(274) xor data_stage(8)(276) xor data_stage(8)(277) xor data_stage(8)(280) xor data_stage(8)(281) xor data_stage(8)(282) xor data_stage(8)(285) xor data_stage(8)(286) xor data_stage(8)(287);
                crc_stage(8)(31) <= crc_stage(7)(31) xor data_stage(8)(256) xor data_stage(8)(259) xor data_stage(8)(263) xor data_stage(8)(268) xor data_stage(8)(274) xor data_stage(8)(277) xor data_stage(8)(281) xor data_stage(8)(283) xor data_stage(8)(284) xor data_stage(8)(285) xor data_stage(8)(287);
            else
                crc_stage(8) <= crc_stage(7);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(9)(39 downto 36) = X"F" then
                crc_stage(9)(0)  <= crc_stage(8)(0) xor data_stage(9)(288) xor data_stage(9)(296) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(311) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(1)  <= crc_stage(8)(1) xor data_stage(9)(289) xor data_stage(9)(297) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(306) xor data_stage(9)(310) xor data_stage(9)(311) xor data_stage(9)(312) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(319);
                crc_stage(9)(2)  <= crc_stage(8)(2) xor data_stage(9)(288) xor data_stage(9)(290) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(306) xor data_stage(9)(307) xor data_stage(9)(311) xor data_stage(9)(312) xor data_stage(9)(313) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(317);
                crc_stage(9)(3)  <= crc_stage(8)(3) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(291) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(305) xor data_stage(9)(306) xor data_stage(9)(307) xor data_stage(9)(308) xor data_stage(9)(312) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(316) xor data_stage(9)(317) xor data_stage(9)(318);
                crc_stage(9)(4)  <= crc_stage(8)(4) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(292) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(307) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(317) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(5)  <= crc_stage(8)(5) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(293) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(6)  <= crc_stage(8)(6) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(294) xor data_stage(9)(296) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(303) xor data_stage(9)(305) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(316) xor data_stage(9)(317) xor data_stage(9)(318);
                crc_stage(9)(7)  <= crc_stage(8)(7) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(295) xor data_stage(9)(297) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(307) xor data_stage(9)(309) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(317) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(8)  <= crc_stage(8)(8) xor data_stage(9)(288) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(296) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(308) xor data_stage(9)(310) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(9)  <= crc_stage(8)(9) xor data_stage(9)(289) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(297) xor data_stage(9)(298) xor data_stage(9)(299) xor data_stage(9)(300) xor data_stage(9)(301) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(310) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(317) xor data_stage(9)(318);
                crc_stage(9)(10) <= crc_stage(8)(10) xor data_stage(9)(288) xor data_stage(9)(290) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(297) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(307) xor data_stage(9)(310) xor data_stage(9)(313) xor data_stage(9)(316) xor data_stage(9)(317);
                crc_stage(9)(11) <= crc_stage(8)(11) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(291) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(308) xor data_stage(9)(311) xor data_stage(9)(314) xor data_stage(9)(317) xor data_stage(9)(318);
                crc_stage(9)(12) <= crc_stage(8)(12) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(292) xor data_stage(9)(296) xor data_stage(9)(297) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(312) xor data_stage(9)(315) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(13) <= crc_stage(8)(13) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(293) xor data_stage(9)(297) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(307) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(313) xor data_stage(9)(316) xor data_stage(9)(319);
                crc_stage(9)(14) <= crc_stage(8)(14) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(294) xor data_stage(9)(298) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(305) xor data_stage(9)(308) xor data_stage(9)(310) xor data_stage(9)(311) xor data_stage(9)(314) xor data_stage(9)(317);
                crc_stage(9)(15) <= crc_stage(8)(15) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(295) xor data_stage(9)(299) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(309) xor data_stage(9)(311) xor data_stage(9)(312) xor data_stage(9)(315) xor data_stage(9)(318);
                crc_stage(9)(16) <= crc_stage(8)(16) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(298) xor data_stage(9)(301) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(307) xor data_stage(9)(309) xor data_stage(9)(311) xor data_stage(9)(312) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(318);
                crc_stage(9)(17) <= crc_stage(8)(17) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(299) xor data_stage(9)(302) xor data_stage(9)(303) xor data_stage(9)(305) xor data_stage(9)(308) xor data_stage(9)(310) xor data_stage(9)(312) xor data_stage(9)(313) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(317) xor data_stage(9)(319);
                crc_stage(9)(18) <= crc_stage(8)(18) xor data_stage(9)(288) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(300) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(309) xor data_stage(9)(311) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(316) xor data_stage(9)(317) xor data_stage(9)(318);
                crc_stage(9)(19) <= crc_stage(8)(19) xor data_stage(9)(289) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(297) xor data_stage(9)(301) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(310) xor data_stage(9)(312) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(317) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(20) <= crc_stage(8)(20) xor data_stage(9)(288) xor data_stage(9)(290) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(297) xor data_stage(9)(300) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(314) xor data_stage(9)(316);
                crc_stage(9)(21) <= crc_stage(8)(21) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(291) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(300) xor data_stage(9)(301) xor data_stage(9)(302) xor data_stage(9)(303) xor data_stage(9)(307) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(317) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(22) <= crc_stage(8)(22) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(292) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(298) xor data_stage(9)(300) xor data_stage(9)(301) xor data_stage(9)(305) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(311) xor data_stage(9)(313);
                crc_stage(9)(23) <= crc_stage(8)(23) xor data_stage(9)(288) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(293) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(302) xor data_stage(9)(306) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(311) xor data_stage(9)(312) xor data_stage(9)(314);
                crc_stage(9)(24) <= crc_stage(8)(24) xor data_stage(9)(288) xor data_stage(9)(289) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(294) xor data_stage(9)(297) xor data_stage(9)(298) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(309) xor data_stage(9)(312) xor data_stage(9)(314) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(25) <= crc_stage(8)(25) xor data_stage(9)(289) xor data_stage(9)(290) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(299) xor data_stage(9)(300) xor data_stage(9)(302) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(311) xor data_stage(9)(314) xor data_stage(9)(318);
                crc_stage(9)(26) <= crc_stage(8)(26) xor data_stage(9)(290) xor data_stage(9)(291) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(296) xor data_stage(9)(297) xor data_stage(9)(300) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(312) xor data_stage(9)(315) xor data_stage(9)(319);
                crc_stage(9)(27) <= crc_stage(8)(27) xor data_stage(9)(291) xor data_stage(9)(292) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(297) xor data_stage(9)(300) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(316) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(28) <= crc_stage(8)(28) xor data_stage(9)(292) xor data_stage(9)(293) xor data_stage(9)(295) xor data_stage(9)(297) xor data_stage(9)(300) xor data_stage(9)(301) xor data_stage(9)(303) xor data_stage(9)(305) xor data_stage(9)(307) xor data_stage(9)(311) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(316) xor data_stage(9)(317) xor data_stage(9)(318);
                crc_stage(9)(29) <= crc_stage(8)(29) xor data_stage(9)(293) xor data_stage(9)(294) xor data_stage(9)(296) xor data_stage(9)(298) xor data_stage(9)(301) xor data_stage(9)(302) xor data_stage(9)(304) xor data_stage(9)(306) xor data_stage(9)(308) xor data_stage(9)(312) xor data_stage(9)(314) xor data_stage(9)(315) xor data_stage(9)(317) xor data_stage(9)(318) xor data_stage(9)(319);
                crc_stage(9)(30) <= crc_stage(8)(30) xor data_stage(9)(294) xor data_stage(9)(295) xor data_stage(9)(296) xor data_stage(9)(297) xor data_stage(9)(298) xor data_stage(9)(299) xor data_stage(9)(300) xor data_stage(9)(304) xor data_stage(9)(307) xor data_stage(9)(310) xor data_stage(9)(311) xor data_stage(9)(314) xor data_stage(9)(316);
                crc_stage(9)(31) <= crc_stage(8)(31) xor data_stage(9)(295) xor data_stage(9)(297) xor data_stage(9)(299) xor data_stage(9)(301) xor data_stage(9)(302) xor data_stage(9)(303) xor data_stage(9)(304) xor data_stage(9)(308) xor data_stage(9)(309) xor data_stage(9)(310) xor data_stage(9)(312) xor data_stage(9)(313) xor data_stage(9)(314) xor data_stage(9)(317) xor data_stage(9)(318) xor data_stage(9)(319);
            else
                crc_stage(9) <= crc_stage(8);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(10)(43 downto 40) = X"F" then
                crc_stage(10)(0)  <= crc_stage(9)(0) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(324) xor data_stage(10)(326) xor data_stage(10)(329) xor data_stage(10)(330) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(345) xor data_stage(10)(346) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(1)  <= crc_stage(9)(1) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(325) xor data_stage(10)(327) xor data_stage(10)(330) xor data_stage(10)(331) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(351);
                crc_stage(10)(2)  <= crc_stage(9)(2) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(331) xor data_stage(10)(332) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(347) xor data_stage(10)(348);
                crc_stage(10)(3)  <= crc_stage(9)(3) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(332) xor data_stage(10)(333) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(346) xor data_stage(10)(348) xor data_stage(10)(349);
                crc_stage(10)(4)  <= crc_stage(9)(4) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(330) xor data_stage(10)(333) xor data_stage(10)(334) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(349) xor data_stage(10)(350);
                crc_stage(10)(5)  <= crc_stage(9)(5) xor data_stage(10)(320) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(331) xor data_stage(10)(334) xor data_stage(10)(335) xor data_stage(10)(345) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(348) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(6)  <= crc_stage(9)(6) xor data_stage(10)(322) xor data_stage(10)(325) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(332) xor data_stage(10)(335) xor data_stage(10)(336) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(345) xor data_stage(10)(347) xor data_stage(10)(348) xor data_stage(10)(349) xor data_stage(10)(350);
                crc_stage(10)(7)  <= crc_stage(9)(7) xor data_stage(10)(323) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(330) xor data_stage(10)(333) xor data_stage(10)(336) xor data_stage(10)(337) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(346) xor data_stage(10)(348) xor data_stage(10)(349) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(8)  <= crc_stage(9)(8) xor data_stage(10)(320) xor data_stage(10)(324) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(330) xor data_stage(10)(331) xor data_stage(10)(334) xor data_stage(10)(337) xor data_stage(10)(338) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(347) xor data_stage(10)(349) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(9)  <= crc_stage(9)(9) xor data_stage(10)(322) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(331) xor data_stage(10)(332) xor data_stage(10)(335) xor data_stage(10)(338) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(344) xor data_stage(10)(348);
                crc_stage(10)(10) <= crc_stage(9)(10) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(327) xor data_stage(10)(332) xor data_stage(10)(333) xor data_stage(10)(336) xor data_stage(10)(339) xor data_stage(10)(346) xor data_stage(10)(349) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(11) <= crc_stage(9)(11) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(333) xor data_stage(10)(334) xor data_stage(10)(337) xor data_stage(10)(340) xor data_stage(10)(347) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(12) <= crc_stage(9)(12) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(334) xor data_stage(10)(335) xor data_stage(10)(338) xor data_stage(10)(341) xor data_stage(10)(348) xor data_stage(10)(351);
                crc_stage(10)(13) <= crc_stage(9)(13) xor data_stage(10)(320) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(330) xor data_stage(10)(335) xor data_stage(10)(336) xor data_stage(10)(339) xor data_stage(10)(342) xor data_stage(10)(349);
                crc_stage(10)(14) <= crc_stage(9)(14) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(331) xor data_stage(10)(336) xor data_stage(10)(337) xor data_stage(10)(340) xor data_stage(10)(343) xor data_stage(10)(350);
                crc_stage(10)(15) <= crc_stage(9)(15) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(330) xor data_stage(10)(332) xor data_stage(10)(337) xor data_stage(10)(338) xor data_stage(10)(341) xor data_stage(10)(344) xor data_stage(10)(351);
                crc_stage(10)(16) <= crc_stage(9)(16) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(331) xor data_stage(10)(333) xor data_stage(10)(338) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(343) xor data_stage(10)(346) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(17) <= crc_stage(9)(17) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(332) xor data_stage(10)(334) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(344) xor data_stage(10)(347) xor data_stage(10)(351);
                crc_stage(10)(18) <= crc_stage(9)(18) xor data_stage(10)(320) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(329) xor data_stage(10)(330) xor data_stage(10)(333) xor data_stage(10)(335) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(345) xor data_stage(10)(348);
                crc_stage(10)(19) <= crc_stage(9)(19) xor data_stage(10)(321) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(330) xor data_stage(10)(331) xor data_stage(10)(334) xor data_stage(10)(336) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(346) xor data_stage(10)(349);
                crc_stage(10)(20) <= crc_stage(9)(20) xor data_stage(10)(321) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(330) xor data_stage(10)(331) xor data_stage(10)(332) xor data_stage(10)(335) xor data_stage(10)(337) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(344) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(351);
                crc_stage(10)(21) <= crc_stage(9)(21) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(324) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(331) xor data_stage(10)(332) xor data_stage(10)(333) xor data_stage(10)(336) xor data_stage(10)(338) xor data_stage(10)(340) xor data_stage(10)(343) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(348) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(22) <= crc_stage(9)(22) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(330) xor data_stage(10)(332) xor data_stage(10)(333) xor data_stage(10)(334) xor data_stage(10)(337) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(348) xor data_stage(10)(349) xor data_stage(10)(350);
                crc_stage(10)(23) <= crc_stage(9)(23) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(331) xor data_stage(10)(333) xor data_stage(10)(334) xor data_stage(10)(335) xor data_stage(10)(338) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(346) xor data_stage(10)(347) xor data_stage(10)(348) xor data_stage(10)(349) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(24) <= crc_stage(9)(24) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(324) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(332) xor data_stage(10)(334) xor data_stage(10)(335) xor data_stage(10)(336) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(347) xor data_stage(10)(348) xor data_stage(10)(349);
                crc_stage(10)(25) <= crc_stage(9)(25) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(328) xor data_stage(10)(333) xor data_stage(10)(335) xor data_stage(10)(336) xor data_stage(10)(337) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(346) xor data_stage(10)(348) xor data_stage(10)(349) xor data_stage(10)(351);
                crc_stage(10)(26) <= crc_stage(9)(26) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(334) xor data_stage(10)(336) xor data_stage(10)(337) xor data_stage(10)(338) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(347) xor data_stage(10)(349) xor data_stage(10)(350);
                crc_stage(10)(27) <= crc_stage(9)(27) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(327) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(335) xor data_stage(10)(337) xor data_stage(10)(338) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(344) xor data_stage(10)(348);
                crc_stage(10)(28) <= crc_stage(9)(28) xor data_stage(10)(321) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(328) xor data_stage(10)(336) xor data_stage(10)(338) xor data_stage(10)(339) xor data_stage(10)(344) xor data_stage(10)(346) xor data_stage(10)(349) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(29) <= crc_stage(9)(29) xor data_stage(10)(322) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(326) xor data_stage(10)(329) xor data_stage(10)(337) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(345) xor data_stage(10)(347) xor data_stage(10)(350) xor data_stage(10)(351);
                crc_stage(10)(30) <= crc_stage(9)(30) xor data_stage(10)(321) xor data_stage(10)(322) xor data_stage(10)(323) xor data_stage(10)(324) xor data_stage(10)(325) xor data_stage(10)(327) xor data_stage(10)(329) xor data_stage(10)(338) xor data_stage(10)(342) xor data_stage(10)(343) xor data_stage(10)(345) xor data_stage(10)(348) xor data_stage(10)(350);
                crc_stage(10)(31) <= crc_stage(9)(31) xor data_stage(10)(320) xor data_stage(10)(321) xor data_stage(10)(323) xor data_stage(10)(325) xor data_stage(10)(328) xor data_stage(10)(329) xor data_stage(10)(339) xor data_stage(10)(340) xor data_stage(10)(341) xor data_stage(10)(342) xor data_stage(10)(344) xor data_stage(10)(345) xor data_stage(10)(349) xor data_stage(10)(350);
            else
                crc_stage(10) <= crc_stage(9);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(11)(47 downto 44) = X"F" then
                crc_stage(11)(0)  <= crc_stage(10)(0) xor data_stage(11)(354) xor data_stage(11)(356) xor data_stage(11)(357) xor data_stage(11)(361) xor data_stage(11)(363) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(380);
                crc_stage(11)(1)  <= crc_stage(10)(1) xor data_stage(11)(352) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(362) xor data_stage(11)(364) xor data_stage(11)(369) xor data_stage(11)(370) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(381);
                crc_stage(11)(2)  <= crc_stage(10)(2) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(356) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(363) xor data_stage(11)(365) xor data_stage(11)(370) xor data_stage(11)(371) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(382);
                crc_stage(11)(3)  <= crc_stage(10)(3) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(357) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(364) xor data_stage(11)(366) xor data_stage(11)(371) xor data_stage(11)(372) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(381) xor data_stage(11)(383);
                crc_stage(11)(4)  <= crc_stage(10)(4) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(358) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(365) xor data_stage(11)(367) xor data_stage(11)(372) xor data_stage(11)(373) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(381) xor data_stage(11)(382);
                crc_stage(11)(5)  <= crc_stage(10)(5) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(359) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(366) xor data_stage(11)(368) xor data_stage(11)(373) xor data_stage(11)(374) xor data_stage(11)(380) xor data_stage(11)(381) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(6)  <= crc_stage(10)(6) xor data_stage(11)(352) xor data_stage(11)(354) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(374) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(380) xor data_stage(11)(381) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(7)  <= crc_stage(10)(7) xor data_stage(11)(353) xor data_stage(11)(355) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(375) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(381) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(8)  <= crc_stage(10)(8) xor data_stage(11)(352) xor data_stage(11)(354) xor data_stage(11)(356) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(364) xor data_stage(11)(369) xor data_stage(11)(370) xor data_stage(11)(376) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(9)  <= crc_stage(10)(9) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(361) xor data_stage(11)(364) xor data_stage(11)(365) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(370) xor data_stage(11)(371) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(381) xor data_stage(11)(383);
                crc_stage(11)(10) <= crc_stage(10)(10) xor data_stage(11)(353) xor data_stage(11)(355) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(365) xor data_stage(11)(366) xor data_stage(11)(368) xor data_stage(11)(370) xor data_stage(11)(371) xor data_stage(11)(372) xor data_stage(11)(375) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(382);
                crc_stage(11)(11) <= crc_stage(10)(11) xor data_stage(11)(352) xor data_stage(11)(354) xor data_stage(11)(356) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(364) xor data_stage(11)(366) xor data_stage(11)(367) xor data_stage(11)(369) xor data_stage(11)(371) xor data_stage(11)(372) xor data_stage(11)(373) xor data_stage(11)(376) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(383);
                crc_stage(11)(12) <= crc_stage(10)(12) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(363) xor data_stage(11)(364) xor data_stage(11)(365) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(370) xor data_stage(11)(372) xor data_stage(11)(373) xor data_stage(11)(374) xor data_stage(11)(377) xor data_stage(11)(380) xor data_stage(11)(381);
                crc_stage(11)(13) <= crc_stage(10)(13) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(356) xor data_stage(11)(358) xor data_stage(11)(364) xor data_stage(11)(365) xor data_stage(11)(366) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(371) xor data_stage(11)(373) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(378) xor data_stage(11)(381) xor data_stage(11)(382);
                crc_stage(11)(14) <= crc_stage(10)(14) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(359) xor data_stage(11)(365) xor data_stage(11)(366) xor data_stage(11)(367) xor data_stage(11)(369) xor data_stage(11)(370) xor data_stage(11)(372) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(379) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(15) <= crc_stage(10)(15) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(358) xor data_stage(11)(360) xor data_stage(11)(366) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(370) xor data_stage(11)(371) xor data_stage(11)(373) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(380) xor data_stage(11)(383);
                crc_stage(11)(16) <= crc_stage(10)(16) xor data_stage(11)(352) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(359) xor data_stage(11)(363) xor data_stage(11)(367) xor data_stage(11)(371) xor data_stage(11)(372) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(380) xor data_stage(11)(381);
                crc_stage(11)(17) <= crc_stage(10)(17) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(360) xor data_stage(11)(364) xor data_stage(11)(368) xor data_stage(11)(372) xor data_stage(11)(373) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(381) xor data_stage(11)(382);
                crc_stage(11)(18) <= crc_stage(10)(18) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(356) xor data_stage(11)(357) xor data_stage(11)(361) xor data_stage(11)(365) xor data_stage(11)(369) xor data_stage(11)(373) xor data_stage(11)(374) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(19) <= crc_stage(10)(19) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(362) xor data_stage(11)(366) xor data_stage(11)(370) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(383);
                crc_stage(11)(20) <= crc_stage(10)(20) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(361) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(371) xor data_stage(11)(377) xor data_stage(11)(379) xor data_stage(11)(380);
                crc_stage(11)(21) <= crc_stage(10)(21) xor data_stage(11)(352) xor data_stage(11)(354) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(370) xor data_stage(11)(372) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(381);
                crc_stage(11)(22) <= crc_stage(10)(22) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(362) xor data_stage(11)(364) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(371) xor data_stage(11)(373) xor data_stage(11)(375) xor data_stage(11)(380) xor data_stage(11)(382);
                crc_stage(11)(23) <= crc_stage(10)(23) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(363) xor data_stage(11)(365) xor data_stage(11)(369) xor data_stage(11)(370) xor data_stage(11)(372) xor data_stage(11)(374) xor data_stage(11)(376) xor data_stage(11)(381) xor data_stage(11)(383);
                crc_stage(11)(24) <= crc_stage(10)(24) xor data_stage(11)(352) xor data_stage(11)(355) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(364) xor data_stage(11)(366) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(370) xor data_stage(11)(371) xor data_stage(11)(373) xor data_stage(11)(376) xor data_stage(11)(378) xor data_stage(11)(380) xor data_stage(11)(382);
                crc_stage(11)(25) <= crc_stage(10)(25) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(357) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(364) xor data_stage(11)(365) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(370) xor data_stage(11)(371) xor data_stage(11)(372) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(381) xor data_stage(11)(383);
                crc_stage(11)(26) <= crc_stage(10)(26) xor data_stage(11)(352) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(358) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(365) xor data_stage(11)(366) xor data_stage(11)(368) xor data_stage(11)(369) xor data_stage(11)(371) xor data_stage(11)(372) xor data_stage(11)(373) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(379) xor data_stage(11)(380) xor data_stage(11)(381) xor data_stage(11)(382);
                crc_stage(11)(27) <= crc_stage(10)(27) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(359) xor data_stage(11)(362) xor data_stage(11)(363) xor data_stage(11)(366) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(370) xor data_stage(11)(372) xor data_stage(11)(373) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(381) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(28) <= crc_stage(10)(28) xor data_stage(11)(355) xor data_stage(11)(357) xor data_stage(11)(358) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(364) xor data_stage(11)(367) xor data_stage(11)(371) xor data_stage(11)(373) xor data_stage(11)(374) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(380) xor data_stage(11)(382) xor data_stage(11)(383);
                crc_stage(11)(29) <= crc_stage(10)(29) xor data_stage(11)(352) xor data_stage(11)(356) xor data_stage(11)(358) xor data_stage(11)(359) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(365) xor data_stage(11)(368) xor data_stage(11)(372) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(381) xor data_stage(11)(383);
                crc_stage(11)(30) <= crc_stage(10)(30) xor data_stage(11)(352) xor data_stage(11)(353) xor data_stage(11)(354) xor data_stage(11)(356) xor data_stage(11)(359) xor data_stage(11)(360) xor data_stage(11)(361) xor data_stage(11)(362) xor data_stage(11)(366) xor data_stage(11)(368) xor data_stage(11)(373) xor data_stage(11)(377) xor data_stage(11)(378) xor data_stage(11)(379) xor data_stage(11)(382);
                crc_stage(11)(31) <= crc_stage(10)(31) xor data_stage(11)(353) xor data_stage(11)(355) xor data_stage(11)(356) xor data_stage(11)(360) xor data_stage(11)(362) xor data_stage(11)(367) xor data_stage(11)(368) xor data_stage(11)(374) xor data_stage(11)(375) xor data_stage(11)(376) xor data_stage(11)(377) xor data_stage(11)(379) xor data_stage(11)(383);
            else
                crc_stage(11) <= crc_stage(10);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(12)(51 downto 48) = X"F" then
                crc_stage(12)(0)  <= crc_stage(11)(0) xor data_stage(12)(384) xor data_stage(12)(385) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(389) xor data_stage(12)(393) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(406) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(411) xor data_stage(12)(413) xor data_stage(12)(414) xor data_stage(12)(415);
                crc_stage(12)(1)  <= crc_stage(11)(1) xor data_stage(12)(385) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(390) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(407) xor data_stage(12)(409) xor data_stage(12)(410) xor data_stage(12)(412) xor data_stage(12)(414) xor data_stage(12)(415);
                crc_stage(12)(2)  <= crc_stage(11)(2) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(391) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(408) xor data_stage(12)(410) xor data_stage(12)(411) xor data_stage(12)(413) xor data_stage(12)(415);
                crc_stage(12)(3)  <= crc_stage(11)(3) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(392) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(409) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(414);
                crc_stage(12)(4)  <= crc_stage(11)(4) xor data_stage(12)(384) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(393) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(410) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(415);
                crc_stage(12)(5)  <= crc_stage(11)(5) xor data_stage(12)(385) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(411) xor data_stage(12)(413) xor data_stage(12)(414);
                crc_stage(12)(6)  <= crc_stage(11)(6) xor data_stage(12)(385) xor data_stage(12)(387) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(396) xor data_stage(12)(398) xor data_stage(12)(400) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(409) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(413);
                crc_stage(12)(7)  <= crc_stage(11)(7) xor data_stage(12)(384) xor data_stage(12)(386) xor data_stage(12)(388) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(395) xor data_stage(12)(397) xor data_stage(12)(399) xor data_stage(12)(401) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(410) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(414);
                crc_stage(12)(8)  <= crc_stage(11)(8) xor data_stage(12)(384) xor data_stage(12)(385) xor data_stage(12)(387) xor data_stage(12)(389) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(394) xor data_stage(12)(396) xor data_stage(12)(398) xor data_stage(12)(400) xor data_stage(12)(402) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(411) xor data_stage(12)(413) xor data_stage(12)(414) xor data_stage(12)(415);
                crc_stage(12)(9)  <= crc_stage(11)(9) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(392) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(410) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(413);
                crc_stage(12)(10) <= crc_stage(11)(10) xor data_stage(12)(385) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(409) xor data_stage(12)(412) xor data_stage(12)(415);
                crc_stage(12)(11) <= crc_stage(11)(11) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(410) xor data_stage(12)(413);
                crc_stage(12)(12) <= crc_stage(11)(12) xor data_stage(12)(384) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(411) xor data_stage(12)(414);
                crc_stage(12)(13) <= crc_stage(11)(13) xor data_stage(12)(385) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(393) xor data_stage(12)(394) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(409) xor data_stage(12)(410) xor data_stage(12)(412) xor data_stage(12)(415);
                crc_stage(12)(14) <= crc_stage(11)(14) xor data_stage(12)(386) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(410) xor data_stage(12)(411) xor data_stage(12)(413);
                crc_stage(12)(15) <= crc_stage(11)(15) xor data_stage(12)(384) xor data_stage(12)(387) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(414);
                crc_stage(12)(16) <= crc_stage(11)(16) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(395) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(403) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(410) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(414);
                crc_stage(12)(17) <= crc_stage(11)(17) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(396) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(404) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(415);
                crc_stage(12)(18) <= crc_stage(11)(18) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(393) xor data_stage(12)(394) xor data_stage(12)(397) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(405) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(414);
                crc_stage(12)(19) <= crc_stage(11)(19) xor data_stage(12)(384) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(398) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(406) xor data_stage(12)(409) xor data_stage(12)(410) xor data_stage(12)(413) xor data_stage(12)(414) xor data_stage(12)(415);
                crc_stage(12)(20) <= crc_stage(11)(20) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(398) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(410) xor data_stage(12)(413);
                crc_stage(12)(21) <= crc_stage(11)(21) xor data_stage(12)(384) xor data_stage(12)(385) xor data_stage(12)(386) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(396) xor data_stage(12)(398) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(410) xor data_stage(12)(413) xor data_stage(12)(415);
                crc_stage(12)(22) <= crc_stage(11)(22) xor data_stage(12)(384) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(394) xor data_stage(12)(396) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(401) xor data_stage(12)(403) xor data_stage(12)(405) xor data_stage(12)(407) xor data_stage(12)(409) xor data_stage(12)(413) xor data_stage(12)(415);
                crc_stage(12)(23) <= crc_stage(11)(23) xor data_stage(12)(385) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(395) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(402) xor data_stage(12)(404) xor data_stage(12)(406) xor data_stage(12)(408) xor data_stage(12)(410) xor data_stage(12)(414);
                crc_stage(12)(24) <= crc_stage(11)(24) xor data_stage(12)(385) xor data_stage(12)(387) xor data_stage(12)(389) xor data_stage(12)(392) xor data_stage(12)(395) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(413) xor data_stage(12)(414);
                crc_stage(12)(25) <= crc_stage(11)(25) xor data_stage(12)(384) xor data_stage(12)(385) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(407) xor data_stage(12)(411) xor data_stage(12)(413);
                crc_stage(12)(26) <= crc_stage(11)(26) xor data_stage(12)(384) xor data_stage(12)(385) xor data_stage(12)(386) xor data_stage(12)(388) xor data_stage(12)(389) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(408) xor data_stage(12)(412) xor data_stage(12)(414);
                crc_stage(12)(27) <= crc_stage(11)(27) xor data_stage(12)(384) xor data_stage(12)(390) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(400) xor data_stage(12)(402) xor data_stage(12)(405) xor data_stage(12)(408) xor data_stage(12)(411) xor data_stage(12)(414);
                crc_stage(12)(28) <= crc_stage(11)(28) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(389) xor data_stage(12)(391) xor data_stage(12)(392) xor data_stage(12)(400) xor data_stage(12)(402) xor data_stage(12)(403) xor data_stage(12)(408) xor data_stage(12)(411) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(414);
                crc_stage(12)(29) <= crc_stage(11)(29) xor data_stage(12)(384) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(390) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(401) xor data_stage(12)(403) xor data_stage(12)(404) xor data_stage(12)(409) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(414) xor data_stage(12)(415);
                crc_stage(12)(30) <= crc_stage(11)(30) xor data_stage(12)(386) xor data_stage(12)(387) xor data_stage(12)(388) xor data_stage(12)(391) xor data_stage(12)(395) xor data_stage(12)(396) xor data_stage(12)(398) xor data_stage(12)(399) xor data_stage(12)(401) xor data_stage(12)(404) xor data_stage(12)(405) xor data_stage(12)(406) xor data_stage(12)(408) xor data_stage(12)(409) xor data_stage(12)(410) xor data_stage(12)(411);
                crc_stage(12)(31) <= crc_stage(11)(31) xor data_stage(12)(384) xor data_stage(12)(385) xor data_stage(12)(386) xor data_stage(12)(388) xor data_stage(12)(392) xor data_stage(12)(393) xor data_stage(12)(394) xor data_stage(12)(395) xor data_stage(12)(397) xor data_stage(12)(398) xor data_stage(12)(400) xor data_stage(12)(401) xor data_stage(12)(405) xor data_stage(12)(407) xor data_stage(12)(408) xor data_stage(12)(410) xor data_stage(12)(412) xor data_stage(12)(413) xor data_stage(12)(414) xor data_stage(12)(415);
            else
                crc_stage(12) <= crc_stage(11);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(13)(55 downto 52) = X"F" then
                crc_stage(13)(0)  <= crc_stage(12)(0) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(425) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(433) xor data_stage(13)(439) xor data_stage(13)(440) xor data_stage(13)(444) xor data_stage(13)(445) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(1)  <= crc_stage(12)(1) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(426) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(434) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(445) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(2)  <= crc_stage(12)(2) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(427) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(435) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(3)  <= crc_stage(12)(3) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(428) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(436) xor data_stage(13)(442) xor data_stage(13)(443) xor data_stage(13)(447);
                crc_stage(13)(4)  <= crc_stage(12)(4) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(429) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(437) xor data_stage(13)(443) xor data_stage(13)(444);
                crc_stage(13)(5)  <= crc_stage(12)(5) xor data_stage(13)(416) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(430) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(438) xor data_stage(13)(444) xor data_stage(13)(445);
                crc_stage(13)(6)  <= crc_stage(12)(6) xor data_stage(13)(416) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(440) xor data_stage(13)(444) xor data_stage(13)(447);
                crc_stage(13)(7)  <= crc_stage(12)(7) xor data_stage(13)(417) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(441) xor data_stage(13)(445);
                crc_stage(13)(8)  <= crc_stage(12)(8) xor data_stage(13)(418) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(439) xor data_stage(13)(442) xor data_stage(13)(446);
                crc_stage(13)(9)  <= crc_stage(12)(9) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(426) xor data_stage(13)(429) xor data_stage(13)(432) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(443) xor data_stage(13)(444) xor data_stage(13)(445) xor data_stage(13)(446);
                crc_stage(13)(10) <= crc_stage(12)(10) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(431) xor data_stage(13)(438) xor data_stage(13)(440);
                crc_stage(13)(11) <= crc_stage(12)(11) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(432) xor data_stage(13)(439) xor data_stage(13)(441);
                crc_stage(13)(12) <= crc_stage(12)(12) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(433) xor data_stage(13)(440) xor data_stage(13)(442);
                crc_stage(13)(13) <= crc_stage(12)(13) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(434) xor data_stage(13)(441) xor data_stage(13)(443);
                crc_stage(13)(14) <= crc_stage(12)(14) xor data_stage(13)(416) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(435) xor data_stage(13)(442) xor data_stage(13)(444);
                crc_stage(13)(15) <= crc_stage(12)(15) xor data_stage(13)(417) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(436) xor data_stage(13)(443) xor data_stage(13)(445);
                crc_stage(13)(16) <= crc_stage(12)(16) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(431) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(437) xor data_stage(13)(439) xor data_stage(13)(440) xor data_stage(13)(445) xor data_stage(13)(447);
                crc_stage(13)(17) <= crc_stage(12)(17) xor data_stage(13)(417) xor data_stage(13)(418) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(432) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(438) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(446);
                crc_stage(13)(18) <= crc_stage(12)(18) xor data_stage(13)(416) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(433) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(439) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(447);
                crc_stage(13)(19) <= crc_stage(12)(19) xor data_stage(13)(417) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(434) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(440) xor data_stage(13)(442) xor data_stage(13)(443);
                crc_stage(13)(20) <= crc_stage(12)(20) xor data_stage(13)(417) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(426) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(433) xor data_stage(13)(435) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(443) xor data_stage(13)(445) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(21) <= crc_stage(12)(21) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(425) xor data_stage(13)(428) xor data_stage(13)(431) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(436) xor data_stage(13)(438) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(445);
                crc_stage(13)(22) <= crc_stage(12)(22) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(437) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(443) xor data_stage(13)(444) xor data_stage(13)(445) xor data_stage(13)(447);
                crc_stage(13)(23) <= crc_stage(12)(23) xor data_stage(13)(416) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(438) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(443) xor data_stage(13)(444) xor data_stage(13)(445) xor data_stage(13)(446);
                crc_stage(13)(24) <= crc_stage(12)(24) xor data_stage(13)(416) xor data_stage(13)(418) xor data_stage(13)(424) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(434) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(440) xor data_stage(13)(442) xor data_stage(13)(443);
                crc_stage(13)(25) <= crc_stage(12)(25) xor data_stage(13)(416) xor data_stage(13)(418) xor data_stage(13)(419) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(435) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(439) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(443) xor data_stage(13)(445) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(26) <= crc_stage(12)(26) xor data_stage(13)(417) xor data_stage(13)(419) xor data_stage(13)(420) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(433) xor data_stage(13)(436) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(439) xor data_stage(13)(440) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(444) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(27) <= crc_stage(12)(27) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(420) xor data_stage(13)(421) xor data_stage(13)(425) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(432) xor data_stage(13)(434) xor data_stage(13)(437) xor data_stage(13)(438) xor data_stage(13)(441) xor data_stage(13)(442) xor data_stage(13)(443) xor data_stage(13)(444) xor data_stage(13)(446);
                crc_stage(13)(28) <= crc_stage(12)(28) xor data_stage(13)(416) xor data_stage(13)(421) xor data_stage(13)(422) xor data_stage(13)(425) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(435) xor data_stage(13)(438) xor data_stage(13)(440) xor data_stage(13)(442) xor data_stage(13)(443) xor data_stage(13)(446);
                crc_stage(13)(29) <= crc_stage(12)(29) xor data_stage(13)(417) xor data_stage(13)(422) xor data_stage(13)(423) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(436) xor data_stage(13)(439) xor data_stage(13)(441) xor data_stage(13)(443) xor data_stage(13)(444) xor data_stage(13)(447);
                crc_stage(13)(30) <= crc_stage(12)(30) xor data_stage(13)(417) xor data_stage(13)(423) xor data_stage(13)(424) xor data_stage(13)(425) xor data_stage(13)(430) xor data_stage(13)(431) xor data_stage(13)(432) xor data_stage(13)(437) xor data_stage(13)(439) xor data_stage(13)(442) xor data_stage(13)(446) xor data_stage(13)(447);
                crc_stage(13)(31) <= crc_stage(12)(31) xor data_stage(13)(416) xor data_stage(13)(417) xor data_stage(13)(424) xor data_stage(13)(426) xor data_stage(13)(427) xor data_stage(13)(428) xor data_stage(13)(429) xor data_stage(13)(430) xor data_stage(13)(432) xor data_stage(13)(438) xor data_stage(13)(439) xor data_stage(13)(443) xor data_stage(13)(444) xor data_stage(13)(445) xor data_stage(13)(446);
            else
                crc_stage(13) <= crc_stage(12);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(14)(59 downto 56) = X"F" then
                crc_stage(14)(0)  <= crc_stage(13)(0) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(454) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(462) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(467) xor data_stage(14)(468) xor data_stage(14)(475) xor data_stage(14)(478);
                crc_stage(14)(1)  <= crc_stage(13)(1) xor data_stage(14)(448) xor data_stage(14)(450) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(455) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(463) xor data_stage(14)(465) xor data_stage(14)(466) xor data_stage(14)(468) xor data_stage(14)(469) xor data_stage(14)(476) xor data_stage(14)(479);
                crc_stage(14)(2)  <= crc_stage(13)(2) xor data_stage(14)(448) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(456) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(464) xor data_stage(14)(466) xor data_stage(14)(467) xor data_stage(14)(469) xor data_stage(14)(470) xor data_stage(14)(477);
                crc_stage(14)(3)  <= crc_stage(13)(3) xor data_stage(14)(448) xor data_stage(14)(449) xor data_stage(14)(450) xor data_stage(14)(452) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(457) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(465) xor data_stage(14)(467) xor data_stage(14)(468) xor data_stage(14)(470) xor data_stage(14)(471) xor data_stage(14)(478);
                crc_stage(14)(4)  <= crc_stage(13)(4) xor data_stage(14)(448) xor data_stage(14)(449) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(458) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(463) xor data_stage(14)(466) xor data_stage(14)(468) xor data_stage(14)(469) xor data_stage(14)(471) xor data_stage(14)(472) xor data_stage(14)(479);
                crc_stage(14)(5)  <= crc_stage(13)(5) xor data_stage(14)(449) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(454) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(459) xor data_stage(14)(462) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(467) xor data_stage(14)(469) xor data_stage(14)(470) xor data_stage(14)(472) xor data_stage(14)(473);
                crc_stage(14)(6)  <= crc_stage(13)(6) xor data_stage(14)(449) xor data_stage(14)(450) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(462) xor data_stage(14)(463) xor data_stage(14)(467) xor data_stage(14)(470) xor data_stage(14)(471) xor data_stage(14)(473) xor data_stage(14)(474) xor data_stage(14)(475) xor data_stage(14)(478);
                crc_stage(14)(7)  <= crc_stage(13)(7) xor data_stage(14)(448) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(468) xor data_stage(14)(471) xor data_stage(14)(472) xor data_stage(14)(474) xor data_stage(14)(475) xor data_stage(14)(476) xor data_stage(14)(479);
                crc_stage(14)(8)  <= crc_stage(13)(8) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(469) xor data_stage(14)(472) xor data_stage(14)(473) xor data_stage(14)(475) xor data_stage(14)(476) xor data_stage(14)(477);
                crc_stage(14)(9)  <= crc_stage(13)(9) xor data_stage(14)(449) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(456) xor data_stage(14)(459) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(466) xor data_stage(14)(467) xor data_stage(14)(468) xor data_stage(14)(470) xor data_stage(14)(473) xor data_stage(14)(474) xor data_stage(14)(475) xor data_stage(14)(476) xor data_stage(14)(477);
                crc_stage(14)(10) <= crc_stage(13)(10) xor data_stage(14)(449) xor data_stage(14)(450) xor data_stage(14)(455) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(462) xor data_stage(14)(469) xor data_stage(14)(471) xor data_stage(14)(474) xor data_stage(14)(476) xor data_stage(14)(477);
                crc_stage(14)(11) <= crc_stage(13)(11) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(456) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(463) xor data_stage(14)(470) xor data_stage(14)(472) xor data_stage(14)(475) xor data_stage(14)(477) xor data_stage(14)(478);
                crc_stage(14)(12) <= crc_stage(13)(12) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(457) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(464) xor data_stage(14)(471) xor data_stage(14)(473) xor data_stage(14)(476) xor data_stage(14)(478) xor data_stage(14)(479);
                crc_stage(14)(13) <= crc_stage(13)(13) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(458) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(463) xor data_stage(14)(465) xor data_stage(14)(472) xor data_stage(14)(474) xor data_stage(14)(477) xor data_stage(14)(479);
                crc_stage(14)(14) <= crc_stage(13)(14) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(459) xor data_stage(14)(462) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(466) xor data_stage(14)(473) xor data_stage(14)(475) xor data_stage(14)(478);
                crc_stage(14)(15) <= crc_stage(13)(15) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(460) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(467) xor data_stage(14)(474) xor data_stage(14)(476) xor data_stage(14)(479);
                crc_stage(14)(16) <= crc_stage(13)(16) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(466) xor data_stage(14)(467) xor data_stage(14)(477) xor data_stage(14)(478);
                crc_stage(14)(17) <= crc_stage(13)(17) xor data_stage(14)(448) xor data_stage(14)(450) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(462) xor data_stage(14)(463) xor data_stage(14)(467) xor data_stage(14)(468) xor data_stage(14)(478) xor data_stage(14)(479);
                crc_stage(14)(18) <= crc_stage(13)(18) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(468) xor data_stage(14)(469) xor data_stage(14)(479);
                crc_stage(14)(19) <= crc_stage(13)(19) xor data_stage(14)(448) xor data_stage(14)(450) xor data_stage(14)(452) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(469) xor data_stage(14)(470);
                crc_stage(14)(20) <= crc_stage(13)(20) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(466) xor data_stage(14)(467) xor data_stage(14)(468) xor data_stage(14)(470) xor data_stage(14)(471) xor data_stage(14)(475) xor data_stage(14)(478);
                crc_stage(14)(21) <= crc_stage(13)(21) xor data_stage(14)(448) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(459) xor data_stage(14)(461) xor data_stage(14)(469) xor data_stage(14)(471) xor data_stage(14)(472) xor data_stage(14)(475) xor data_stage(14)(476) xor data_stage(14)(478) xor data_stage(14)(479);
                crc_stage(14)(22) <= crc_stage(13)(22) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(456) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(467) xor data_stage(14)(468) xor data_stage(14)(470) xor data_stage(14)(472) xor data_stage(14)(473) xor data_stage(14)(475) xor data_stage(14)(476) xor data_stage(14)(477) xor data_stage(14)(478) xor data_stage(14)(479);
                crc_stage(14)(23) <= crc_stage(13)(23) xor data_stage(14)(448) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(454) xor data_stage(14)(457) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(465) xor data_stage(14)(466) xor data_stage(14)(468) xor data_stage(14)(469) xor data_stage(14)(471) xor data_stage(14)(473) xor data_stage(14)(474) xor data_stage(14)(476) xor data_stage(14)(477) xor data_stage(14)(478) xor data_stage(14)(479);
                crc_stage(14)(24) <= crc_stage(13)(24) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(455) xor data_stage(14)(457) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(466) xor data_stage(14)(468) xor data_stage(14)(469) xor data_stage(14)(470) xor data_stage(14)(472) xor data_stage(14)(474) xor data_stage(14)(477) xor data_stage(14)(479);
                crc_stage(14)(25) <= crc_stage(13)(25) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(455) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(464) xor data_stage(14)(466) xor data_stage(14)(468) xor data_stage(14)(469) xor data_stage(14)(470) xor data_stage(14)(471) xor data_stage(14)(473);
                crc_stage(14)(26) <= crc_stage(13)(26) xor data_stage(14)(448) xor data_stage(14)(450) xor data_stage(14)(452) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(465) xor data_stage(14)(467) xor data_stage(14)(469) xor data_stage(14)(470) xor data_stage(14)(471) xor data_stage(14)(472) xor data_stage(14)(474);
                crc_stage(14)(27) <= crc_stage(13)(27) xor data_stage(14)(448) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(461) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(466) xor data_stage(14)(467) xor data_stage(14)(470) xor data_stage(14)(471) xor data_stage(14)(472) xor data_stage(14)(473) xor data_stage(14)(478);
                crc_stage(14)(28) <= crc_stage(13)(28) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(455) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(466) xor data_stage(14)(471) xor data_stage(14)(472) xor data_stage(14)(473) xor data_stage(14)(474) xor data_stage(14)(475) xor data_stage(14)(478) xor data_stage(14)(479);
                crc_stage(14)(29) <= crc_stage(13)(29) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(454) xor data_stage(14)(456) xor data_stage(14)(458) xor data_stage(14)(459) xor data_stage(14)(460) xor data_stage(14)(467) xor data_stage(14)(472) xor data_stage(14)(473) xor data_stage(14)(474) xor data_stage(14)(475) xor data_stage(14)(476) xor data_stage(14)(479);
                crc_stage(14)(30) <= crc_stage(13)(30) xor data_stage(14)(448) xor data_stage(14)(449) xor data_stage(14)(451) xor data_stage(14)(452) xor data_stage(14)(453) xor data_stage(14)(455) xor data_stage(14)(458) xor data_stage(14)(460) xor data_stage(14)(461) xor data_stage(14)(462) xor data_stage(14)(464) xor data_stage(14)(465) xor data_stage(14)(467) xor data_stage(14)(473) xor data_stage(14)(474) xor data_stage(14)(476) xor data_stage(14)(477) xor data_stage(14)(478);
                crc_stage(14)(31) <= crc_stage(13)(31) xor data_stage(14)(448) xor data_stage(14)(450) xor data_stage(14)(451) xor data_stage(14)(453) xor data_stage(14)(456) xor data_stage(14)(457) xor data_stage(14)(458) xor data_stage(14)(461) xor data_stage(14)(463) xor data_stage(14)(464) xor data_stage(14)(466) xor data_stage(14)(467) xor data_stage(14)(474) xor data_stage(14)(477) xor data_stage(14)(479);
            else
                crc_stage(14) <= crc_stage(13);
            end if;
        end if;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if keep_stage(15)(63 downto 60) = X"F" then
                crc_stage(15)(0)  <= crc_stage(14)(0) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(26) xor crcIn(29) xor crcIn(30) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(481) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(496) xor data_stage(15)(500) xor data_stage(15)(502) xor data_stage(15)(503) xor data_stage(15)(506);
                crc_stage(15)(1)  <= crc_stage(14)(1) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor crcIn(30) xor crcIn(31) xor data_stage(15)(481) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(489) xor data_stage(15)(497) xor data_stage(15)(501) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(507);
                crc_stage(15)(2)  <= crc_stage(14)(2) xor crcIn(0) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(6) xor crcIn(7) xor crcIn(8) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(28) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(488) xor data_stage(15)(489) xor data_stage(15)(490) xor data_stage(15)(498) xor data_stage(15)(502) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(508);
                crc_stage(15)(3)  <= crc_stage(14)(3) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(7) xor crcIn(8) xor crcIn(9) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(29) xor data_stage(15)(481) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(489) xor data_stage(15)(490) xor data_stage(15)(491) xor data_stage(15)(499) xor data_stage(15)(503) xor data_stage(15)(505) xor data_stage(15)(506) xor data_stage(15)(509);
                crc_stage(15)(4)  <= crc_stage(14)(4) xor crcIn(0) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(10) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(28) xor crcIn(30) xor data_stage(15)(482) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(490) xor data_stage(15)(491) xor data_stage(15)(492) xor data_stage(15)(500) xor data_stage(15)(504) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(510);
                crc_stage(15)(5)  <= crc_stage(14)(5) xor crcIn(1) xor crcIn(3) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(11) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(28) xor crcIn(29) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(483) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(489) xor data_stage(15)(491) xor data_stage(15)(492) xor data_stage(15)(493) xor data_stage(15)(501) xor data_stage(15)(505) xor data_stage(15)(507) xor data_stage(15)(508) xor data_stage(15)(511);
                crc_stage(15)(6)  <= crc_stage(14)(6) xor crcIn(1) xor crcIn(5) xor crcIn(7) xor crcIn(8) xor crcIn(16) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(25) xor crcIn(27) xor crcIn(28) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(489) xor data_stage(15)(490) xor data_stage(15)(492) xor data_stage(15)(493) xor data_stage(15)(494) xor data_stage(15)(496) xor data_stage(15)(500) xor data_stage(15)(503) xor data_stage(15)(508) xor data_stage(15)(509);
                crc_stage(15)(7)  <= crc_stage(14)(7) xor crcIn(0) xor crcIn(2) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(17) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(26) xor crcIn(28) xor crcIn(29) xor data_stage(15)(481) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(490) xor data_stage(15)(491) xor data_stage(15)(493) xor data_stage(15)(494) xor data_stage(15)(495) xor data_stage(15)(497) xor data_stage(15)(501) xor data_stage(15)(504) xor data_stage(15)(509) xor data_stage(15)(510);
                crc_stage(15)(8)  <= crc_stage(14)(8) xor crcIn(0) xor crcIn(1) xor crcIn(3) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(18) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(27) xor crcIn(29) xor crcIn(30) xor data_stage(15)(480) xor data_stage(15)(482) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(491) xor data_stage(15)(492) xor data_stage(15)(494) xor data_stage(15)(495) xor data_stage(15)(496) xor data_stage(15)(498) xor data_stage(15)(502) xor data_stage(15)(505) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(9)  <= crc_stage(14)(9) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(12) xor crcIn(17) xor crcIn(18) xor crcIn(20) xor crcIn(21) xor crcIn(25) xor crcIn(26) xor crcIn(28) xor crcIn(29) xor data_stage(15)(480) xor data_stage(15)(482) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(492) xor data_stage(15)(493) xor data_stage(15)(495) xor data_stage(15)(497) xor data_stage(15)(499) xor data_stage(15)(500) xor data_stage(15)(502) xor data_stage(15)(511);
                crc_stage(15)(10) <= crc_stage(14)(10) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(17) xor crcIn(20) xor crcIn(23) xor crcIn(24) xor crcIn(27) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(482) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(487) xor data_stage(15)(489) xor data_stage(15)(493) xor data_stage(15)(494) xor data_stage(15)(498) xor data_stage(15)(501) xor data_stage(15)(502) xor data_stage(15)(506);
                crc_stage(15)(11) <= crc_stage(14)(11) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(18) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(28) xor data_stage(15)(481) xor data_stage(15)(483) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(488) xor data_stage(15)(490) xor data_stage(15)(494) xor data_stage(15)(495) xor data_stage(15)(499) xor data_stage(15)(502) xor data_stage(15)(503) xor data_stage(15)(507);
                crc_stage(15)(12) <= crc_stage(14)(12) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(6) xor crcIn(7) xor crcIn(9) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(19) xor crcIn(22) xor crcIn(25) xor crcIn(26) xor crcIn(29) xor data_stage(15)(482) xor data_stage(15)(484) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(489) xor data_stage(15)(491) xor data_stage(15)(495) xor data_stage(15)(496) xor data_stage(15)(500) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(508);
                crc_stage(15)(13) <= crc_stage(14)(13) xor crcIn(0) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(7) xor crcIn(8) xor crcIn(10) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(20) xor crcIn(23) xor crcIn(26) xor crcIn(27) xor crcIn(30) xor data_stage(15)(480) xor data_stage(15)(483) xor data_stage(15)(485) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(490) xor data_stage(15)(492) xor data_stage(15)(496) xor data_stage(15)(497) xor data_stage(15)(501) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(509);
                crc_stage(15)(14) <= crc_stage(14)(14) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(11) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(21) xor crcIn(24) xor crcIn(27) xor crcIn(28) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(481) xor data_stage(15)(484) xor data_stage(15)(486) xor data_stage(15)(488) xor data_stage(15)(489) xor data_stage(15)(491) xor data_stage(15)(493) xor data_stage(15)(497) xor data_stage(15)(498) xor data_stage(15)(502) xor data_stage(15)(505) xor data_stage(15)(506) xor data_stage(15)(510);
                crc_stage(15)(15) <= crc_stage(14)(15) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(12) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(22) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor data_stage(15)(481) xor data_stage(15)(482) xor data_stage(15)(485) xor data_stage(15)(487) xor data_stage(15)(489) xor data_stage(15)(490) xor data_stage(15)(492) xor data_stage(15)(494) xor data_stage(15)(498) xor data_stage(15)(499) xor data_stage(15)(503) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(511);
                crc_stage(15)(16) <= crc_stage(14)(16) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(7) xor crcIn(8) xor crcIn(12) xor crcIn(13) xor crcIn(15) xor crcIn(16) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(24) xor crcIn(31) xor data_stage(15)(481) xor data_stage(15)(484) xor data_stage(15)(487) xor data_stage(15)(490) xor data_stage(15)(491) xor data_stage(15)(493) xor data_stage(15)(495) xor data_stage(15)(496) xor data_stage(15)(499) xor data_stage(15)(502) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(508);
                crc_stage(15)(17) <= crc_stage(14)(17) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(8) xor crcIn(9) xor crcIn(13) xor crcIn(14) xor crcIn(16) xor crcIn(17) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(25) xor data_stage(15)(482) xor data_stage(15)(485) xor data_stage(15)(488) xor data_stage(15)(491) xor data_stage(15)(492) xor data_stage(15)(494) xor data_stage(15)(496) xor data_stage(15)(497) xor data_stage(15)(500) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(507) xor data_stage(15)(508) xor data_stage(15)(509);
                crc_stage(15)(18) <= crc_stage(14)(18) xor crcIn(0) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(9) xor crcIn(10) xor crcIn(14) xor crcIn(15) xor crcIn(17) xor crcIn(18) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(26) xor data_stage(15)(480) xor data_stage(15)(483) xor data_stage(15)(486) xor data_stage(15)(489) xor data_stage(15)(492) xor data_stage(15)(493) xor data_stage(15)(495) xor data_stage(15)(497) xor data_stage(15)(498) xor data_stage(15)(501) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(506) xor data_stage(15)(508) xor data_stage(15)(509) xor data_stage(15)(510);
                crc_stage(15)(19) <= crc_stage(14)(19) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(10) xor crcIn(11) xor crcIn(15) xor crcIn(16) xor crcIn(18) xor crcIn(19) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor data_stage(15)(480) xor data_stage(15)(481) xor data_stage(15)(484) xor data_stage(15)(487) xor data_stage(15)(490) xor data_stage(15)(493) xor data_stage(15)(494) xor data_stage(15)(496) xor data_stage(15)(498) xor data_stage(15)(499) xor data_stage(15)(502) xor data_stage(15)(505) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(509) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(20) <= crc_stage(14)(20) xor crcIn(0) xor crcIn(1) xor crcIn(7) xor crcIn(8) xor crcIn(10) xor crcIn(16) xor crcIn(18) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor crcIn(30) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(491) xor data_stage(15)(494) xor data_stage(15)(495) xor data_stage(15)(496) xor data_stage(15)(497) xor data_stage(15)(499) xor data_stage(15)(502) xor data_stage(15)(507) xor data_stage(15)(508) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(21) <= crc_stage(14)(21) xor crcIn(0) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(10) xor crcIn(12) xor crcIn(18) xor crcIn(20) xor crcIn(21) xor data_stage(15)(480) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(485) xor data_stage(15)(492) xor data_stage(15)(495) xor data_stage(15)(497) xor data_stage(15)(498) xor data_stage(15)(502) xor data_stage(15)(506) xor data_stage(15)(508) xor data_stage(15)(509) xor data_stage(15)(511);
                crc_stage(15)(22) <= crc_stage(14)(22) xor crcIn(2) xor crcIn(4) xor crcIn(7) xor crcIn(9) xor crcIn(12) xor crcIn(13) xor crcIn(17) xor crcIn(18) xor crcIn(20) xor crcIn(23) xor crcIn(24) xor crcIn(26) xor crcIn(29) xor crcIn(30) xor crcIn(31) xor data_stage(15)(482) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(493) xor data_stage(15)(498) xor data_stage(15)(499) xor data_stage(15)(500) xor data_stage(15)(502) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(509) xor data_stage(15)(510);
                crc_stage(15)(23) <= crc_stage(14)(23) xor crcIn(3) xor crcIn(5) xor crcIn(8) xor crcIn(10) xor crcIn(13) xor crcIn(14) xor crcIn(18) xor crcIn(19) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor crcIn(30) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(483) xor data_stage(15)(488) xor data_stage(15)(489) xor data_stage(15)(494) xor data_stage(15)(499) xor data_stage(15)(500) xor data_stage(15)(501) xor data_stage(15)(503) xor data_stage(15)(507) xor data_stage(15)(508) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(24) <= crc_stage(14)(24) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(5) xor crcIn(9) xor crcIn(10) xor crcIn(12) xor crcIn(14) xor crcIn(15) xor crcIn(17) xor crcIn(18) xor crcIn(21) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor crcIn(30) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(488) xor data_stage(15)(489) xor data_stage(15)(490) xor data_stage(15)(495) xor data_stage(15)(496) xor data_stage(15)(501) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(506) xor data_stage(15)(508) xor data_stage(15)(509) xor data_stage(15)(511);
                crc_stage(15)(25) <= crc_stage(14)(25) xor crcIn(0) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(12) xor crcIn(13) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(20) xor crcIn(21) xor crcIn(23) xor crcIn(25) xor data_stage(15)(481) xor data_stage(15)(482) xor data_stage(15)(486) xor data_stage(15)(489) xor data_stage(15)(490) xor data_stage(15)(491) xor data_stage(15)(497) xor data_stage(15)(500) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(509) xor data_stage(15)(510);
                crc_stage(15)(26) <= crc_stage(14)(26) xor crcIn(0) xor crcIn(1) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(13) xor crcIn(14) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(21) xor crcIn(22) xor crcIn(24) xor crcIn(26) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(487) xor data_stage(15)(490) xor data_stage(15)(491) xor data_stage(15)(492) xor data_stage(15)(498) xor data_stage(15)(501) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(506) xor data_stage(15)(507) xor data_stage(15)(508) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(27) <= crc_stage(14)(27) xor crcIn(0) xor crcIn(4) xor crcIn(7) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(14) xor crcIn(15) xor crcIn(20) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(29) xor crcIn(30) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(481) xor data_stage(15)(482) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(491) xor data_stage(15)(492) xor data_stage(15)(493) xor data_stage(15)(496) xor data_stage(15)(499) xor data_stage(15)(500) xor data_stage(15)(503) xor data_stage(15)(505) xor data_stage(15)(507) xor data_stage(15)(508) xor data_stage(15)(509) xor data_stage(15)(511);
                crc_stage(15)(28) <= crc_stage(14)(28) xor crcIn(2) xor crcIn(4) xor crcIn(6) xor crcIn(8) xor crcIn(10) xor crcIn(13) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor crcIn(28) xor crcIn(29) xor data_stage(15)(480) xor data_stage(15)(484) xor data_stage(15)(486) xor data_stage(15)(492) xor data_stage(15)(493) xor data_stage(15)(494) xor data_stage(15)(496) xor data_stage(15)(497) xor data_stage(15)(501) xor data_stage(15)(502) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(508) xor data_stage(15)(509) xor data_stage(15)(510);
                crc_stage(15)(29) <= crc_stage(14)(29) xor crcIn(3) xor crcIn(5) xor crcIn(7) xor crcIn(9) xor crcIn(11) xor crcIn(14) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(28) xor crcIn(29) xor crcIn(30) xor data_stage(15)(480) xor data_stage(15)(481) xor data_stage(15)(485) xor data_stage(15)(487) xor data_stage(15)(493) xor data_stage(15)(494) xor data_stage(15)(495) xor data_stage(15)(497) xor data_stage(15)(498) xor data_stage(15)(502) xor data_stage(15)(503) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(509) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(30) <= crc_stage(14)(30) xor crcIn(1) xor crcIn(2) xor crcIn(5) xor crcIn(8) xor crcIn(11) xor crcIn(15) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor data_stage(15)(483) xor data_stage(15)(484) xor data_stage(15)(487) xor data_stage(15)(494) xor data_stage(15)(495) xor data_stage(15)(498) xor data_stage(15)(499) xor data_stage(15)(500) xor data_stage(15)(502) xor data_stage(15)(504) xor data_stage(15)(505) xor data_stage(15)(510) xor data_stage(15)(511);
                crc_stage(15)(31) <= crc_stage(14)(31) xor crcIn(0) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(9) xor crcIn(10) xor crcIn(11) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor crcIn(30) xor crcIn(31) xor data_stage(15)(480) xor data_stage(15)(481) xor data_stage(15)(482) xor data_stage(15)(483) xor data_stage(15)(485) xor data_stage(15)(486) xor data_stage(15)(487) xor data_stage(15)(495) xor data_stage(15)(499) xor data_stage(15)(501) xor data_stage(15)(502) xor data_stage(15)(505) xor data_stage(15)(511);
            else
                crc_stage(15)(0)  <= crc_stage(14)(0) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(26) xor crcIn(29) xor crcIn(30) xor crcIn(31);
                crc_stage(15)(1)  <= crc_stage(14)(1) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor crcIn(30) xor crcIn(31);
                crc_stage(15)(2)  <= crc_stage(14)(2) xor crcIn(0) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(6) xor crcIn(7) xor crcIn(8) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(28) xor crcIn(31);
                crc_stage(15)(3)  <= crc_stage(14)(3) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(7) xor crcIn(8) xor crcIn(9) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(29);
                crc_stage(15)(4)  <= crc_stage(14)(4) xor crcIn(0) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(10) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(28);
                crc_stage(15)(5)  <= crc_stage(14)(5) xor crcIn(1) xor crcIn(3) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(11) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(28) xor crcIn(29) xor crcIn(31);
                crc_stage(15)(6)  <= crc_stage(14)(6) xor crcIn(1) xor crcIn(5) xor crcIn(7) xor crcIn(8) xor crcIn(16) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(25) xor crcIn(27) xor crcIn(28) xor crcIn(31);
                crc_stage(15)(7)  <= crc_stage(14)(7) xor crcIn(0) xor crcIn(2) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(17) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(26) xor crcIn(28) xor crcIn(29);
                crc_stage(15)(8)  <= crc_stage(14)(8) xor crcIn(0) xor crcIn(1) xor crcIn(3) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(18) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(27) xor crcIn(29) xor crcIn(30);
                crc_stage(15)(9)  <= crc_stage(14)(9) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(12) xor crcIn(17) xor crcIn(18) xor crcIn(20) xor crcIn(21) xor crcIn(25) xor crcIn(26) xor crcIn(28) xor crcIn(29);
                crc_stage(15)(10) <= crc_stage(14)(10) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(17) xor crcIn(20) xor crcIn(23) xor crcIn(24) xor crcIn(27) xor crcIn(31);
                crc_stage(15)(11) <= crc_stage(14)(11) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(18) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(28);
                crc_stage(15)(12) <= crc_stage(14)(12) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(6) xor crcIn(7) xor crcIn(9) xor crcIn(11) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(19) xor crcIn(22) xor crcIn(25) xor crcIn(26) xor crcIn(29);
                crc_stage(15)(13) <= crc_stage(14)(13) xor crcIn(0) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(7) xor crcIn(8) xor crcIn(10) xor crcIn(12) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(20) xor crcIn(23) xor crcIn(26) xor crcIn(27) xor crcIn(30);
                crc_stage(15)(14) <= crc_stage(14)(14) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(11) xor crcIn(13) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(21) xor crcIn(24) xor crcIn(27) xor crcIn(28) xor crcIn(31);
                crc_stage(15)(15) <= crc_stage(14)(15) xor crcIn(2) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(9) xor crcIn(10) xor crcIn(12) xor crcIn(14) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(22) xor crcIn(25) xor crcIn(28) xor crcIn(29);
                crc_stage(15)(16) <= crc_stage(14)(16) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(7) xor crcIn(8) xor crcIn(12) xor crcIn(13) xor crcIn(15) xor crcIn(16) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(24) xor crcIn(31);
                crc_stage(15)(17) <= crc_stage(14)(17) xor crcIn(1) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(8) xor crcIn(9) xor crcIn(13) xor crcIn(14) xor crcIn(16) xor crcIn(17) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(25);
                crc_stage(15)(18) <= crc_stage(14)(18) xor crcIn(0) xor crcIn(2) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(9) xor crcIn(10) xor crcIn(14) xor crcIn(15) xor crcIn(17) xor crcIn(18) xor crcIn(22) xor crcIn(23) xor crcIn(24) xor crcIn(26);
                crc_stage(15)(19) <= crc_stage(14)(19) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(7) xor crcIn(10) xor crcIn(11) xor crcIn(15) xor crcIn(16) xor crcIn(18) xor crcIn(19) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27);
                crc_stage(15)(20) <= crc_stage(14)(20) xor crcIn(0) xor crcIn(1) xor crcIn(7) xor crcIn(8) xor crcIn(10) xor crcIn(16) xor crcIn(18) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor crcIn(30) xor crcIn(31);
                crc_stage(15)(21) <= crc_stage(14)(21) xor crcIn(0) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(8) xor crcIn(9) xor crcIn(10) xor crcIn(12) xor crcIn(18) xor crcIn(20) xor crcIn(21);
                crc_stage(15)(22) <= crc_stage(14)(22) xor crcIn(2) xor crcIn(4) xor crcIn(7) xor crcIn(9) xor crcIn(12) xor crcIn(13) xor crcIn(17) xor crcIn(18) xor crcIn(20) xor crcIn(23) xor crcIn(24) xor crcIn(26) xor crcIn(29) xor crcIn(30) xor crcIn(31);
                crc_stage(15)(23) <= crc_stage(14)(23) xor crcIn(3) xor crcIn(5) xor crcIn(8) xor crcIn(10) xor crcIn(13) xor crcIn(14) xor crcIn(18) xor crcIn(19) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor crcIn(30) xor crcIn(31);
                crc_stage(15)(24) <= crc_stage(14)(24) xor crcIn(0) xor crcIn(1) xor crcIn(2) xor crcIn(5) xor crcIn(9) xor crcIn(10) xor crcIn(12) xor crcIn(14) xor crcIn(15) xor crcIn(17) xor crcIn(18) xor crcIn(21) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor crcIn(30);
                crc_stage(15)(25) <= crc_stage(14)(25) xor crcIn(0) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(12) xor crcIn(13) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(20) xor crcIn(21) xor crcIn(23) xor crcIn(25);
                crc_stage(15)(26) <= crc_stage(14)(26) xor crcIn(0) xor crcIn(1) xor crcIn(4) xor crcIn(5) xor crcIn(6) xor crcIn(13) xor crcIn(14) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(21) xor crcIn(22) xor crcIn(24) xor crcIn(26);
                crc_stage(15)(27) <= crc_stage(14)(27) xor crcIn(0) xor crcIn(4) xor crcIn(7) xor crcIn(10) xor crcIn(11) xor crcIn(12) xor crcIn(14) xor crcIn(15) xor crcIn(20) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(27) xor crcIn(29) xor crcIn(30) xor crcIn(31);
                crc_stage(15)(28) <= crc_stage(14)(28) xor crcIn(2) xor crcIn(4) xor crcIn(6) xor crcIn(8) xor crcIn(10) xor crcIn(13) xor crcIn(15) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27) xor crcIn(28) xor crcIn(29);
                crc_stage(15)(29) <= crc_stage(14)(29) xor crcIn(3) xor crcIn(5) xor crcIn(7) xor crcIn(9) xor crcIn(11) xor crcIn(14) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(24) xor crcIn(25) xor crcIn(26) xor crcIn(28) xor crcIn(29) xor crcIn(30);
                crc_stage(15)(30) <= crc_stage(14)(30) xor crcIn(1) xor crcIn(2) xor crcIn(5) xor crcIn(8) xor crcIn(11) xor crcIn(15) xor crcIn(23) xor crcIn(24) xor crcIn(25) xor crcIn(27);
                crc_stage(15)(31) <= crc_stage(14)(31) xor crcIn(0) xor crcIn(1) xor crcIn(3) xor crcIn(4) xor crcIn(5) xor crcIn(9) xor crcIn(10) xor crcIn(11) xor crcIn(16) xor crcIn(17) xor crcIn(18) xor crcIn(19) xor crcIn(20) xor crcIn(21) xor crcIn(22) xor crcIn(23) xor crcIn(25) xor crcIn(28) xor crcIn(29) xor crcIn(30) xor crcIn(31);
            end if;
        end if;
    end process;

    reverse_out_g : if REVERSE_RESULT generate
        reverse_g : for i in 0 to 31 generate
            crcOut(i) <= crc_stage(7)(31 - i) xor FINXOR(31 - i);
        end generate;
    else generate
        crcOut <= crc_stage(7) xor FINXOR;
    end generate;

    reverse_deb_g : for i in 0 to 31 generate
        crc_rev(i) <= crc_stage(7)(31 - i) xor FINXOR(31 - i);
    end generate;

    valid_crc_out <= valid_shreg(valid_shreg'high);

end architecture Behavioral;
