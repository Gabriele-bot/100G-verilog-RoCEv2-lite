`timescale 1ns / 1ps

package Board_params;

    parameter RoCE_CLOCK_PERIOD = 1000/280.00142; // in ns
    parameter MAC_CLOCK_PERIOD = 1000/391; // in ns

    parameter RoCE_DATA_WIDTH = 2048;
  
endpackage
